library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"ff87eb49",
     1 => x"78c848d0",
     2 => x"731e4f26",
     3 => x"c24b711e",
     4 => x"02bfe4f6",
     5 => x"ebc287c3",
     6 => x"48d0ff87",
     7 => x"7378c9c8",
     8 => x"b1e0c049",
     9 => x"7148d4ff",
    10 => x"d8f6c278",
    11 => x"c878c048",
    12 => x"87c50266",
    13 => x"c249ffc3",
    14 => x"c249c087",
    15 => x"cc59e0f6",
    16 => x"87c60266",
    17 => x"4ad5d5c5",
    18 => x"ffcf87c4",
    19 => x"f6c24aff",
    20 => x"f6c25ae4",
    21 => x"78c148e4",
    22 => x"4d2687c4",
    23 => x"4b264c26",
    24 => x"5e0e4f26",
    25 => x"0e5d5c5b",
    26 => x"f6c24a71",
    27 => x"724cbfe0",
    28 => x"87cb029a",
    29 => x"c291c849",
    30 => x"714bc0c0",
    31 => x"c287c483",
    32 => x"c04bc0c4",
    33 => x"7449134d",
    34 => x"dcf6c299",
    35 => x"d4ffb9bf",
    36 => x"c1787148",
    37 => x"c8852cb7",
    38 => x"e804adb7",
    39 => x"d8f6c287",
    40 => x"80c848bf",
    41 => x"58dcf6c2",
    42 => x"1e87effe",
    43 => x"4b711e73",
    44 => x"029a4a13",
    45 => x"497287cb",
    46 => x"1387e7fe",
    47 => x"f5059a4a",
    48 => x"87dafe87",
    49 => x"d8f6c21e",
    50 => x"f6c249bf",
    51 => x"a1c148d8",
    52 => x"b7c0c478",
    53 => x"87db03a9",
    54 => x"c248d4ff",
    55 => x"78bfdcf6",
    56 => x"bfd8f6c2",
    57 => x"d8f6c249",
    58 => x"78a1c148",
    59 => x"a9b7c0c4",
    60 => x"ff87e504",
    61 => x"78c848d0",
    62 => x"48e4f6c2",
    63 => x"4f2678c0",
    64 => x"00000000",
    65 => x"00000000",
    66 => x"5f000000",
    67 => x"0000005f",
    68 => x"00030300",
    69 => x"00000303",
    70 => x"147f7f14",
    71 => x"00147f7f",
    72 => x"6b2e2400",
    73 => x"00123a6b",
    74 => x"18366a4c",
    75 => x"0032566c",
    76 => x"594f7e30",
    77 => x"40683a77",
    78 => x"07040000",
    79 => x"00000003",
    80 => x"3e1c0000",
    81 => x"00004163",
    82 => x"63410000",
    83 => x"00001c3e",
    84 => x"1c3e2a08",
    85 => x"082a3e1c",
    86 => x"3e080800",
    87 => x"0008083e",
    88 => x"e0800000",
    89 => x"00000060",
    90 => x"08080800",
    91 => x"00080808",
    92 => x"60000000",
    93 => x"00000060",
    94 => x"18306040",
    95 => x"0103060c",
    96 => x"597f3e00",
    97 => x"003e7f4d",
    98 => x"7f060400",
    99 => x"0000007f",
   100 => x"71634200",
   101 => x"00464f59",
   102 => x"49632200",
   103 => x"00367f49",
   104 => x"13161c18",
   105 => x"00107f7f",
   106 => x"45672700",
   107 => x"00397d45",
   108 => x"4b7e3c00",
   109 => x"00307949",
   110 => x"71010100",
   111 => x"00070f79",
   112 => x"497f3600",
   113 => x"00367f49",
   114 => x"494f0600",
   115 => x"001e3f69",
   116 => x"66000000",
   117 => x"00000066",
   118 => x"e6800000",
   119 => x"00000066",
   120 => x"14080800",
   121 => x"00222214",
   122 => x"14141400",
   123 => x"00141414",
   124 => x"14222200",
   125 => x"00080814",
   126 => x"51030200",
   127 => x"00060f59",
   128 => x"5d417f3e",
   129 => x"001e1f55",
   130 => x"097f7e00",
   131 => x"007e7f09",
   132 => x"497f7f00",
   133 => x"00367f49",
   134 => x"633e1c00",
   135 => x"00414141",
   136 => x"417f7f00",
   137 => x"001c3e63",
   138 => x"497f7f00",
   139 => x"00414149",
   140 => x"097f7f00",
   141 => x"00010109",
   142 => x"417f3e00",
   143 => x"007a7b49",
   144 => x"087f7f00",
   145 => x"007f7f08",
   146 => x"7f410000",
   147 => x"0000417f",
   148 => x"40602000",
   149 => x"003f7f40",
   150 => x"1c087f7f",
   151 => x"00416336",
   152 => x"407f7f00",
   153 => x"00404040",
   154 => x"0c067f7f",
   155 => x"007f7f06",
   156 => x"0c067f7f",
   157 => x"007f7f18",
   158 => x"417f3e00",
   159 => x"003e7f41",
   160 => x"097f7f00",
   161 => x"00060f09",
   162 => x"61417f3e",
   163 => x"00407e7f",
   164 => x"097f7f00",
   165 => x"00667f19",
   166 => x"4d6f2600",
   167 => x"00327b59",
   168 => x"7f010100",
   169 => x"0001017f",
   170 => x"407f3f00",
   171 => x"003f7f40",
   172 => x"703f0f00",
   173 => x"000f3f70",
   174 => x"18307f7f",
   175 => x"007f7f30",
   176 => x"1c366341",
   177 => x"4163361c",
   178 => x"7c060301",
   179 => x"0103067c",
   180 => x"4d597161",
   181 => x"00414347",
   182 => x"7f7f0000",
   183 => x"00004141",
   184 => x"0c060301",
   185 => x"40603018",
   186 => x"41410000",
   187 => x"00007f7f",
   188 => x"03060c08",
   189 => x"00080c06",
   190 => x"80808080",
   191 => x"00808080",
   192 => x"03000000",
   193 => x"00000407",
   194 => x"54742000",
   195 => x"00787c54",
   196 => x"447f7f00",
   197 => x"00387c44",
   198 => x"447c3800",
   199 => x"00004444",
   200 => x"447c3800",
   201 => x"007f7f44",
   202 => x"547c3800",
   203 => x"00185c54",
   204 => x"7f7e0400",
   205 => x"00000505",
   206 => x"a4bc1800",
   207 => x"007cfca4",
   208 => x"047f7f00",
   209 => x"00787c04",
   210 => x"3d000000",
   211 => x"0000407d",
   212 => x"80808000",
   213 => x"00007dfd",
   214 => x"107f7f00",
   215 => x"00446c38",
   216 => x"3f000000",
   217 => x"0000407f",
   218 => x"180c7c7c",
   219 => x"00787c0c",
   220 => x"047c7c00",
   221 => x"00787c04",
   222 => x"447c3800",
   223 => x"00387c44",
   224 => x"24fcfc00",
   225 => x"00183c24",
   226 => x"243c1800",
   227 => x"00fcfc24",
   228 => x"047c7c00",
   229 => x"00080c04",
   230 => x"545c4800",
   231 => x"00207454",
   232 => x"7f3f0400",
   233 => x"00004444",
   234 => x"407c3c00",
   235 => x"007c7c40",
   236 => x"603c1c00",
   237 => x"001c3c60",
   238 => x"30607c3c",
   239 => x"003c7c60",
   240 => x"10386c44",
   241 => x"00446c38",
   242 => x"e0bc1c00",
   243 => x"001c3c60",
   244 => x"74644400",
   245 => x"00444c5c",
   246 => x"3e080800",
   247 => x"00414177",
   248 => x"7f000000",
   249 => x"0000007f",
   250 => x"77414100",
   251 => x"0008083e",
   252 => x"03010102",
   253 => x"00010202",
   254 => x"7f7f7f7f",
   255 => x"007f7f7f",
   256 => x"1c1c0808",
   257 => x"7f7f3e3e",
   258 => x"3e3e7f7f",
   259 => x"08081c1c",
   260 => x"7c181000",
   261 => x"0010187c",
   262 => x"7c301000",
   263 => x"0010307c",
   264 => x"60603010",
   265 => x"00061e78",
   266 => x"183c6642",
   267 => x"0042663c",
   268 => x"c26a3878",
   269 => x"00386cc6",
   270 => x"60000060",
   271 => x"00600000",
   272 => x"5c5b5e0e",
   273 => x"711e0e5d",
   274 => x"f5f6c24c",
   275 => x"4bc04dbf",
   276 => x"ab741ec0",
   277 => x"c487c702",
   278 => x"78c048a6",
   279 => x"a6c487c5",
   280 => x"c478c148",
   281 => x"49731e66",
   282 => x"c887dfee",
   283 => x"49e0c086",
   284 => x"c487efef",
   285 => x"496a4aa5",
   286 => x"f187f0f0",
   287 => x"85cb87c6",
   288 => x"b7c883c1",
   289 => x"c7ff04ab",
   290 => x"4d262687",
   291 => x"4b264c26",
   292 => x"711e4f26",
   293 => x"f9f6c24a",
   294 => x"f9f6c25a",
   295 => x"4978c748",
   296 => x"2687ddfe",
   297 => x"1e731e4f",
   298 => x"b7c04a71",
   299 => x"87d303aa",
   300 => x"bfc5e0c2",
   301 => x"c187c405",
   302 => x"c087c24b",
   303 => x"c9e0c24b",
   304 => x"c287c45b",
   305 => x"c25ac9e0",
   306 => x"4abfc5e0",
   307 => x"c0c19ac1",
   308 => x"e8ec49a2",
   309 => x"c248fc87",
   310 => x"78bfc5e0",
   311 => x"1e87effe",
   312 => x"66c44a71",
   313 => x"ff49721e",
   314 => x"2687e9df",
   315 => x"c21e4f26",
   316 => x"49bfc5e0",
   317 => x"87d9dcff",
   318 => x"48edf6c2",
   319 => x"c278bfe8",
   320 => x"ec48e9f6",
   321 => x"f6c278bf",
   322 => x"494abfed",
   323 => x"c899ffc3",
   324 => x"48722ab7",
   325 => x"f6c2b071",
   326 => x"4f2658f5",
   327 => x"5c5b5e0e",
   328 => x"4b710e5d",
   329 => x"c287c7ff",
   330 => x"c048e8f6",
   331 => x"ff497350",
   332 => x"7087fedb",
   333 => x"9cc24c49",
   334 => x"cb49eecb",
   335 => x"497087cf",
   336 => x"e8f6c24d",
   337 => x"c105bf97",
   338 => x"66d087e4",
   339 => x"f1f6c249",
   340 => x"d70599bf",
   341 => x"4966d487",
   342 => x"bfe9f6c2",
   343 => x"87cc0599",
   344 => x"dbff4973",
   345 => x"987087cb",
   346 => x"87c2c102",
   347 => x"fdfd4cc1",
   348 => x"ca497587",
   349 => x"987087e3",
   350 => x"c287c602",
   351 => x"c148e8f6",
   352 => x"e8f6c250",
   353 => x"c005bf97",
   354 => x"f6c287e4",
   355 => x"d049bff1",
   356 => x"ff059966",
   357 => x"f6c287d6",
   358 => x"d449bfe9",
   359 => x"ff059966",
   360 => x"497387ca",
   361 => x"87c9daff",
   362 => x"fe059870",
   363 => x"487487fe",
   364 => x"0e87d7fb",
   365 => x"5d5c5b5e",
   366 => x"c086f40e",
   367 => x"bfec4c4d",
   368 => x"48a6c47e",
   369 => x"bff5f6c2",
   370 => x"c01ec178",
   371 => x"fd49c71e",
   372 => x"86c887ca",
   373 => x"ce029870",
   374 => x"fb49ff87",
   375 => x"dac187c7",
   376 => x"ccd9ff49",
   377 => x"c24dc187",
   378 => x"bf97e8f6",
   379 => x"c987c302",
   380 => x"f6c287c0",
   381 => x"c24bbfed",
   382 => x"05bfc5e0",
   383 => x"c387ebc0",
   384 => x"d8ff49fd",
   385 => x"fac387eb",
   386 => x"e4d8ff49",
   387 => x"c3497387",
   388 => x"1e7199ff",
   389 => x"c6fb49c0",
   390 => x"c8497387",
   391 => x"1e7129b7",
   392 => x"fafa49c1",
   393 => x"c686c887",
   394 => x"f6c287c1",
   395 => x"9b4bbff1",
   396 => x"c287dd02",
   397 => x"49bfc1e0",
   398 => x"7087dec7",
   399 => x"87c40598",
   400 => x"87d24bc0",
   401 => x"c749e0c2",
   402 => x"e0c287c3",
   403 => x"87c658c5",
   404 => x"48c1e0c2",
   405 => x"497378c0",
   406 => x"ce0599c2",
   407 => x"49ebc387",
   408 => x"87cdd7ff",
   409 => x"99c24970",
   410 => x"fb87c202",
   411 => x"c149734c",
   412 => x"87ce0599",
   413 => x"ff49f4c3",
   414 => x"7087f6d6",
   415 => x"0299c249",
   416 => x"4cfa87c2",
   417 => x"99c84973",
   418 => x"c387ce05",
   419 => x"d6ff49f5",
   420 => x"497087df",
   421 => x"d50299c2",
   422 => x"f9f6c287",
   423 => x"87ca02bf",
   424 => x"c288c148",
   425 => x"c058fdf6",
   426 => x"4cff87c2",
   427 => x"49734dc1",
   428 => x"ce0599c4",
   429 => x"49f2c387",
   430 => x"87f5d5ff",
   431 => x"99c24970",
   432 => x"c287dc02",
   433 => x"7ebff9f6",
   434 => x"a8b7c748",
   435 => x"87cbc003",
   436 => x"80c1486e",
   437 => x"58fdf6c2",
   438 => x"fe87c2c0",
   439 => x"c34dc14c",
   440 => x"d5ff49fd",
   441 => x"497087cb",
   442 => x"c00299c2",
   443 => x"f6c287d5",
   444 => x"c002bff9",
   445 => x"f6c287c9",
   446 => x"78c048f9",
   447 => x"fd87c2c0",
   448 => x"c34dc14c",
   449 => x"d4ff49fa",
   450 => x"497087e7",
   451 => x"c00299c2",
   452 => x"f6c287d9",
   453 => x"c748bff9",
   454 => x"c003a8b7",
   455 => x"f6c287c9",
   456 => x"78c748f9",
   457 => x"fc87c2c0",
   458 => x"c04dc14c",
   459 => x"c003acb7",
   460 => x"66c487d1",
   461 => x"82d8c14a",
   462 => x"c6c0026a",
   463 => x"744b6a87",
   464 => x"c00f7349",
   465 => x"1ef0c31e",
   466 => x"f749dac1",
   467 => x"86c887ce",
   468 => x"c0029870",
   469 => x"a6c887e2",
   470 => x"f9f6c248",
   471 => x"66c878bf",
   472 => x"c491cb49",
   473 => x"80714866",
   474 => x"bf6e7e70",
   475 => x"87c8c002",
   476 => x"c84bbf6e",
   477 => x"0f734966",
   478 => x"c0029d75",
   479 => x"f6c287c8",
   480 => x"f249bff9",
   481 => x"e0c287fa",
   482 => x"c002bfc9",
   483 => x"c24987dd",
   484 => x"987087c7",
   485 => x"87d3c002",
   486 => x"bff9f6c2",
   487 => x"87e0f249",
   488 => x"c0f449c0",
   489 => x"c9e0c287",
   490 => x"f478c048",
   491 => x"87daf38e",
   492 => x"5c5b5e0e",
   493 => x"711e0e5d",
   494 => x"f5f6c24c",
   495 => x"cdc149bf",
   496 => x"d1c14da1",
   497 => x"747e6981",
   498 => x"87cf029c",
   499 => x"744ba5c4",
   500 => x"f5f6c27b",
   501 => x"f9f249bf",
   502 => x"747b6e87",
   503 => x"87c4059c",
   504 => x"87c24bc0",
   505 => x"49734bc1",
   506 => x"d487faf2",
   507 => x"87c70266",
   508 => x"7087da49",
   509 => x"c087c24a",
   510 => x"cde0c24a",
   511 => x"c9f2265a",
   512 => x"00000087",
   513 => x"00000000",
   514 => x"00000000",
   515 => x"4a711e00",
   516 => x"49bfc8ff",
   517 => x"2648a172",
   518 => x"c8ff1e4f",
   519 => x"c0fe89bf",
   520 => x"c0c0c0c0",
   521 => x"87c401a9",
   522 => x"87c24ac0",
   523 => x"48724ac1",
   524 => x"c21e4f26",
   525 => x"49bfdbe1",
   526 => x"e1c2b9c1",
   527 => x"d4ff59df",
   528 => x"78ffc348",
   529 => x"c048d0ff",
   530 => x"d4ff78e1",
   531 => x"c478c148",
   532 => x"ff787131",
   533 => x"e0c048d0",
   534 => x"004f2678",
   535 => x"0e000000",
   536 => x"5d5c5b5e",
   537 => x"e9f6c20e",
   538 => x"e3c24abf",
   539 => x"4c49bfc8",
   540 => x"4d71bc72",
   541 => x"87e0c7ff",
   542 => x"49744bc0",
   543 => x"c00299d0",
   544 => x"d0ff87e7",
   545 => x"78e1c848",
   546 => x"c548d4ff",
   547 => x"d0497578",
   548 => x"87c30299",
   549 => x"c278f0c3",
   550 => x"7349f6e3",
   551 => x"ff481181",
   552 => x"ff7808d4",
   553 => x"e0c048d0",
   554 => x"2d2cc178",
   555 => x"04abc883",
   556 => x"ff87c7ff",
   557 => x"c287d9c6",
   558 => x"c248c8e3",
   559 => x"78bfe9f6",
   560 => x"4c264d26",
   561 => x"4f264b26",
   562 => x"00000000",
   563 => x"c3e7c11e",
   564 => x"c250de48",
   565 => x"fe49dfe3",
   566 => x"c087eada",
   567 => x"504f2648",
   568 => x"4d4b4355",
   569 => x"41317e41",
   570 => x"1e004352",
   571 => x"fd87c4f3",
   572 => x"87f887ed",
   573 => x"1e164f26",
   574 => x"362e2526",
   575 => x"362e3e3d",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
