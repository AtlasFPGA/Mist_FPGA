
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"ff",x"87",x"eb",x"49"),
     1 => (x"78",x"c8",x"48",x"d0"),
     2 => (x"73",x"1e",x"4f",x"26"),
     3 => (x"c2",x"4b",x"71",x"1e"),
     4 => (x"02",x"bf",x"e4",x"f6"),
     5 => (x"eb",x"c2",x"87",x"c3"),
     6 => (x"48",x"d0",x"ff",x"87"),
     7 => (x"73",x"78",x"c9",x"c8"),
     8 => (x"b1",x"e0",x"c0",x"49"),
     9 => (x"71",x"48",x"d4",x"ff"),
    10 => (x"d8",x"f6",x"c2",x"78"),
    11 => (x"c8",x"78",x"c0",x"48"),
    12 => (x"87",x"c5",x"02",x"66"),
    13 => (x"c2",x"49",x"ff",x"c3"),
    14 => (x"c2",x"49",x"c0",x"87"),
    15 => (x"cc",x"59",x"e0",x"f6"),
    16 => (x"87",x"c6",x"02",x"66"),
    17 => (x"4a",x"d5",x"d5",x"c5"),
    18 => (x"ff",x"cf",x"87",x"c4"),
    19 => (x"f6",x"c2",x"4a",x"ff"),
    20 => (x"f6",x"c2",x"5a",x"e4"),
    21 => (x"78",x"c1",x"48",x"e4"),
    22 => (x"4d",x"26",x"87",x"c4"),
    23 => (x"4b",x"26",x"4c",x"26"),
    24 => (x"5e",x"0e",x"4f",x"26"),
    25 => (x"0e",x"5d",x"5c",x"5b"),
    26 => (x"f6",x"c2",x"4a",x"71"),
    27 => (x"72",x"4c",x"bf",x"e0"),
    28 => (x"87",x"cb",x"02",x"9a"),
    29 => (x"c2",x"91",x"c8",x"49"),
    30 => (x"71",x"4b",x"c0",x"c0"),
    31 => (x"c2",x"87",x"c4",x"83"),
    32 => (x"c0",x"4b",x"c0",x"c4"),
    33 => (x"74",x"49",x"13",x"4d"),
    34 => (x"dc",x"f6",x"c2",x"99"),
    35 => (x"d4",x"ff",x"b9",x"bf"),
    36 => (x"c1",x"78",x"71",x"48"),
    37 => (x"c8",x"85",x"2c",x"b7"),
    38 => (x"e8",x"04",x"ad",x"b7"),
    39 => (x"d8",x"f6",x"c2",x"87"),
    40 => (x"80",x"c8",x"48",x"bf"),
    41 => (x"58",x"dc",x"f6",x"c2"),
    42 => (x"1e",x"87",x"ef",x"fe"),
    43 => (x"4b",x"71",x"1e",x"73"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cb"),
    46 => (x"13",x"87",x"e7",x"fe"),
    47 => (x"f5",x"05",x"9a",x"4a"),
    48 => (x"87",x"da",x"fe",x"87"),
    49 => (x"d8",x"f6",x"c2",x"1e"),
    50 => (x"f6",x"c2",x"49",x"bf"),
    51 => (x"a1",x"c1",x"48",x"d8"),
    52 => (x"b7",x"c0",x"c4",x"78"),
    53 => (x"87",x"db",x"03",x"a9"),
    54 => (x"c2",x"48",x"d4",x"ff"),
    55 => (x"78",x"bf",x"dc",x"f6"),
    56 => (x"bf",x"d8",x"f6",x"c2"),
    57 => (x"d8",x"f6",x"c2",x"49"),
    58 => (x"78",x"a1",x"c1",x"48"),
    59 => (x"a9",x"b7",x"c0",x"c4"),
    60 => (x"ff",x"87",x"e5",x"04"),
    61 => (x"78",x"c8",x"48",x"d0"),
    62 => (x"48",x"e4",x"f6",x"c2"),
    63 => (x"4f",x"26",x"78",x"c0"),
    64 => (x"00",x"00",x"00",x"00"),
    65 => (x"00",x"00",x"00",x"00"),
    66 => (x"5f",x"00",x"00",x"00"),
    67 => (x"00",x"00",x"00",x"5f"),
    68 => (x"00",x"03",x"03",x"00"),
    69 => (x"00",x"00",x"03",x"03"),
    70 => (x"14",x"7f",x"7f",x"14"),
    71 => (x"00",x"14",x"7f",x"7f"),
    72 => (x"6b",x"2e",x"24",x"00"),
    73 => (x"00",x"12",x"3a",x"6b"),
    74 => (x"18",x"36",x"6a",x"4c"),
    75 => (x"00",x"32",x"56",x"6c"),
    76 => (x"59",x"4f",x"7e",x"30"),
    77 => (x"40",x"68",x"3a",x"77"),
    78 => (x"07",x"04",x"00",x"00"),
    79 => (x"00",x"00",x"00",x"03"),
    80 => (x"3e",x"1c",x"00",x"00"),
    81 => (x"00",x"00",x"41",x"63"),
    82 => (x"63",x"41",x"00",x"00"),
    83 => (x"00",x"00",x"1c",x"3e"),
    84 => (x"1c",x"3e",x"2a",x"08"),
    85 => (x"08",x"2a",x"3e",x"1c"),
    86 => (x"3e",x"08",x"08",x"00"),
    87 => (x"00",x"08",x"08",x"3e"),
    88 => (x"e0",x"80",x"00",x"00"),
    89 => (x"00",x"00",x"00",x"60"),
    90 => (x"08",x"08",x"08",x"00"),
    91 => (x"00",x"08",x"08",x"08"),
    92 => (x"60",x"00",x"00",x"00"),
    93 => (x"00",x"00",x"00",x"60"),
    94 => (x"18",x"30",x"60",x"40"),
    95 => (x"01",x"03",x"06",x"0c"),
    96 => (x"59",x"7f",x"3e",x"00"),
    97 => (x"00",x"3e",x"7f",x"4d"),
    98 => (x"7f",x"06",x"04",x"00"),
    99 => (x"00",x"00",x"00",x"7f"),
   100 => (x"71",x"63",x"42",x"00"),
   101 => (x"00",x"46",x"4f",x"59"),
   102 => (x"49",x"63",x"22",x"00"),
   103 => (x"00",x"36",x"7f",x"49"),
   104 => (x"13",x"16",x"1c",x"18"),
   105 => (x"00",x"10",x"7f",x"7f"),
   106 => (x"45",x"67",x"27",x"00"),
   107 => (x"00",x"39",x"7d",x"45"),
   108 => (x"4b",x"7e",x"3c",x"00"),
   109 => (x"00",x"30",x"79",x"49"),
   110 => (x"71",x"01",x"01",x"00"),
   111 => (x"00",x"07",x"0f",x"79"),
   112 => (x"49",x"7f",x"36",x"00"),
   113 => (x"00",x"36",x"7f",x"49"),
   114 => (x"49",x"4f",x"06",x"00"),
   115 => (x"00",x"1e",x"3f",x"69"),
   116 => (x"66",x"00",x"00",x"00"),
   117 => (x"00",x"00",x"00",x"66"),
   118 => (x"e6",x"80",x"00",x"00"),
   119 => (x"00",x"00",x"00",x"66"),
   120 => (x"14",x"08",x"08",x"00"),
   121 => (x"00",x"22",x"22",x"14"),
   122 => (x"14",x"14",x"14",x"00"),
   123 => (x"00",x"14",x"14",x"14"),
   124 => (x"14",x"22",x"22",x"00"),
   125 => (x"00",x"08",x"08",x"14"),
   126 => (x"51",x"03",x"02",x"00"),
   127 => (x"00",x"06",x"0f",x"59"),
   128 => (x"5d",x"41",x"7f",x"3e"),
   129 => (x"00",x"1e",x"1f",x"55"),
   130 => (x"09",x"7f",x"7e",x"00"),
   131 => (x"00",x"7e",x"7f",x"09"),
   132 => (x"49",x"7f",x"7f",x"00"),
   133 => (x"00",x"36",x"7f",x"49"),
   134 => (x"63",x"3e",x"1c",x"00"),
   135 => (x"00",x"41",x"41",x"41"),
   136 => (x"41",x"7f",x"7f",x"00"),
   137 => (x"00",x"1c",x"3e",x"63"),
   138 => (x"49",x"7f",x"7f",x"00"),
   139 => (x"00",x"41",x"41",x"49"),
   140 => (x"09",x"7f",x"7f",x"00"),
   141 => (x"00",x"01",x"01",x"09"),
   142 => (x"41",x"7f",x"3e",x"00"),
   143 => (x"00",x"7a",x"7b",x"49"),
   144 => (x"08",x"7f",x"7f",x"00"),
   145 => (x"00",x"7f",x"7f",x"08"),
   146 => (x"7f",x"41",x"00",x"00"),
   147 => (x"00",x"00",x"41",x"7f"),
   148 => (x"40",x"60",x"20",x"00"),
   149 => (x"00",x"3f",x"7f",x"40"),
   150 => (x"1c",x"08",x"7f",x"7f"),
   151 => (x"00",x"41",x"63",x"36"),
   152 => (x"40",x"7f",x"7f",x"00"),
   153 => (x"00",x"40",x"40",x"40"),
   154 => (x"0c",x"06",x"7f",x"7f"),
   155 => (x"00",x"7f",x"7f",x"06"),
   156 => (x"0c",x"06",x"7f",x"7f"),
   157 => (x"00",x"7f",x"7f",x"18"),
   158 => (x"41",x"7f",x"3e",x"00"),
   159 => (x"00",x"3e",x"7f",x"41"),
   160 => (x"09",x"7f",x"7f",x"00"),
   161 => (x"00",x"06",x"0f",x"09"),
   162 => (x"61",x"41",x"7f",x"3e"),
   163 => (x"00",x"40",x"7e",x"7f"),
   164 => (x"09",x"7f",x"7f",x"00"),
   165 => (x"00",x"66",x"7f",x"19"),
   166 => (x"4d",x"6f",x"26",x"00"),
   167 => (x"00",x"32",x"7b",x"59"),
   168 => (x"7f",x"01",x"01",x"00"),
   169 => (x"00",x"01",x"01",x"7f"),
   170 => (x"40",x"7f",x"3f",x"00"),
   171 => (x"00",x"3f",x"7f",x"40"),
   172 => (x"70",x"3f",x"0f",x"00"),
   173 => (x"00",x"0f",x"3f",x"70"),
   174 => (x"18",x"30",x"7f",x"7f"),
   175 => (x"00",x"7f",x"7f",x"30"),
   176 => (x"1c",x"36",x"63",x"41"),
   177 => (x"41",x"63",x"36",x"1c"),
   178 => (x"7c",x"06",x"03",x"01"),
   179 => (x"01",x"03",x"06",x"7c"),
   180 => (x"4d",x"59",x"71",x"61"),
   181 => (x"00",x"41",x"43",x"47"),
   182 => (x"7f",x"7f",x"00",x"00"),
   183 => (x"00",x"00",x"41",x"41"),
   184 => (x"0c",x"06",x"03",x"01"),
   185 => (x"40",x"60",x"30",x"18"),
   186 => (x"41",x"41",x"00",x"00"),
   187 => (x"00",x"00",x"7f",x"7f"),
   188 => (x"03",x"06",x"0c",x"08"),
   189 => (x"00",x"08",x"0c",x"06"),
   190 => (x"80",x"80",x"80",x"80"),
   191 => (x"00",x"80",x"80",x"80"),
   192 => (x"03",x"00",x"00",x"00"),
   193 => (x"00",x"00",x"04",x"07"),
   194 => (x"54",x"74",x"20",x"00"),
   195 => (x"00",x"78",x"7c",x"54"),
   196 => (x"44",x"7f",x"7f",x"00"),
   197 => (x"00",x"38",x"7c",x"44"),
   198 => (x"44",x"7c",x"38",x"00"),
   199 => (x"00",x"00",x"44",x"44"),
   200 => (x"44",x"7c",x"38",x"00"),
   201 => (x"00",x"7f",x"7f",x"44"),
   202 => (x"54",x"7c",x"38",x"00"),
   203 => (x"00",x"18",x"5c",x"54"),
   204 => (x"7f",x"7e",x"04",x"00"),
   205 => (x"00",x"00",x"05",x"05"),
   206 => (x"a4",x"bc",x"18",x"00"),
   207 => (x"00",x"7c",x"fc",x"a4"),
   208 => (x"04",x"7f",x"7f",x"00"),
   209 => (x"00",x"78",x"7c",x"04"),
   210 => (x"3d",x"00",x"00",x"00"),
   211 => (x"00",x"00",x"40",x"7d"),
   212 => (x"80",x"80",x"80",x"00"),
   213 => (x"00",x"00",x"7d",x"fd"),
   214 => (x"10",x"7f",x"7f",x"00"),
   215 => (x"00",x"44",x"6c",x"38"),
   216 => (x"3f",x"00",x"00",x"00"),
   217 => (x"00",x"00",x"40",x"7f"),
   218 => (x"18",x"0c",x"7c",x"7c"),
   219 => (x"00",x"78",x"7c",x"0c"),
   220 => (x"04",x"7c",x"7c",x"00"),
   221 => (x"00",x"78",x"7c",x"04"),
   222 => (x"44",x"7c",x"38",x"00"),
   223 => (x"00",x"38",x"7c",x"44"),
   224 => (x"24",x"fc",x"fc",x"00"),
   225 => (x"00",x"18",x"3c",x"24"),
   226 => (x"24",x"3c",x"18",x"00"),
   227 => (x"00",x"fc",x"fc",x"24"),
   228 => (x"04",x"7c",x"7c",x"00"),
   229 => (x"00",x"08",x"0c",x"04"),
   230 => (x"54",x"5c",x"48",x"00"),
   231 => (x"00",x"20",x"74",x"54"),
   232 => (x"7f",x"3f",x"04",x"00"),
   233 => (x"00",x"00",x"44",x"44"),
   234 => (x"40",x"7c",x"3c",x"00"),
   235 => (x"00",x"7c",x"7c",x"40"),
   236 => (x"60",x"3c",x"1c",x"00"),
   237 => (x"00",x"1c",x"3c",x"60"),
   238 => (x"30",x"60",x"7c",x"3c"),
   239 => (x"00",x"3c",x"7c",x"60"),
   240 => (x"10",x"38",x"6c",x"44"),
   241 => (x"00",x"44",x"6c",x"38"),
   242 => (x"e0",x"bc",x"1c",x"00"),
   243 => (x"00",x"1c",x"3c",x"60"),
   244 => (x"74",x"64",x"44",x"00"),
   245 => (x"00",x"44",x"4c",x"5c"),
   246 => (x"3e",x"08",x"08",x"00"),
   247 => (x"00",x"41",x"41",x"77"),
   248 => (x"7f",x"00",x"00",x"00"),
   249 => (x"00",x"00",x"00",x"7f"),
   250 => (x"77",x"41",x"41",x"00"),
   251 => (x"00",x"08",x"08",x"3e"),
   252 => (x"03",x"01",x"01",x"02"),
   253 => (x"00",x"01",x"02",x"02"),
   254 => (x"7f",x"7f",x"7f",x"7f"),
   255 => (x"00",x"7f",x"7f",x"7f"),
   256 => (x"1c",x"1c",x"08",x"08"),
   257 => (x"7f",x"7f",x"3e",x"3e"),
   258 => (x"3e",x"3e",x"7f",x"7f"),
   259 => (x"08",x"08",x"1c",x"1c"),
   260 => (x"7c",x"18",x"10",x"00"),
   261 => (x"00",x"10",x"18",x"7c"),
   262 => (x"7c",x"30",x"10",x"00"),
   263 => (x"00",x"10",x"30",x"7c"),
   264 => (x"60",x"60",x"30",x"10"),
   265 => (x"00",x"06",x"1e",x"78"),
   266 => (x"18",x"3c",x"66",x"42"),
   267 => (x"00",x"42",x"66",x"3c"),
   268 => (x"c2",x"6a",x"38",x"78"),
   269 => (x"00",x"38",x"6c",x"c6"),
   270 => (x"60",x"00",x"00",x"60"),
   271 => (x"00",x"60",x"00",x"00"),
   272 => (x"5c",x"5b",x"5e",x"0e"),
   273 => (x"71",x"1e",x"0e",x"5d"),
   274 => (x"f5",x"f6",x"c2",x"4c"),
   275 => (x"4b",x"c0",x"4d",x"bf"),
   276 => (x"ab",x"74",x"1e",x"c0"),
   277 => (x"c4",x"87",x"c7",x"02"),
   278 => (x"78",x"c0",x"48",x"a6"),
   279 => (x"a6",x"c4",x"87",x"c5"),
   280 => (x"c4",x"78",x"c1",x"48"),
   281 => (x"49",x"73",x"1e",x"66"),
   282 => (x"c8",x"87",x"df",x"ee"),
   283 => (x"49",x"e0",x"c0",x"86"),
   284 => (x"c4",x"87",x"ef",x"ef"),
   285 => (x"49",x"6a",x"4a",x"a5"),
   286 => (x"f1",x"87",x"f0",x"f0"),
   287 => (x"85",x"cb",x"87",x"c6"),
   288 => (x"b7",x"c8",x"83",x"c1"),
   289 => (x"c7",x"ff",x"04",x"ab"),
   290 => (x"4d",x"26",x"26",x"87"),
   291 => (x"4b",x"26",x"4c",x"26"),
   292 => (x"71",x"1e",x"4f",x"26"),
   293 => (x"f9",x"f6",x"c2",x"4a"),
   294 => (x"f9",x"f6",x"c2",x"5a"),
   295 => (x"49",x"78",x"c7",x"48"),
   296 => (x"26",x"87",x"dd",x"fe"),
   297 => (x"1e",x"73",x"1e",x"4f"),
   298 => (x"b7",x"c0",x"4a",x"71"),
   299 => (x"87",x"d3",x"03",x"aa"),
   300 => (x"bf",x"c5",x"e0",x"c2"),
   301 => (x"c1",x"87",x"c4",x"05"),
   302 => (x"c0",x"87",x"c2",x"4b"),
   303 => (x"c9",x"e0",x"c2",x"4b"),
   304 => (x"c2",x"87",x"c4",x"5b"),
   305 => (x"c2",x"5a",x"c9",x"e0"),
   306 => (x"4a",x"bf",x"c5",x"e0"),
   307 => (x"c0",x"c1",x"9a",x"c1"),
   308 => (x"e8",x"ec",x"49",x"a2"),
   309 => (x"c2",x"48",x"fc",x"87"),
   310 => (x"78",x"bf",x"c5",x"e0"),
   311 => (x"1e",x"87",x"ef",x"fe"),
   312 => (x"66",x"c4",x"4a",x"71"),
   313 => (x"ff",x"49",x"72",x"1e"),
   314 => (x"26",x"87",x"e9",x"df"),
   315 => (x"c2",x"1e",x"4f",x"26"),
   316 => (x"49",x"bf",x"c5",x"e0"),
   317 => (x"87",x"d9",x"dc",x"ff"),
   318 => (x"48",x"ed",x"f6",x"c2"),
   319 => (x"c2",x"78",x"bf",x"e8"),
   320 => (x"ec",x"48",x"e9",x"f6"),
   321 => (x"f6",x"c2",x"78",x"bf"),
   322 => (x"49",x"4a",x"bf",x"ed"),
   323 => (x"c8",x"99",x"ff",x"c3"),
   324 => (x"48",x"72",x"2a",x"b7"),
   325 => (x"f6",x"c2",x"b0",x"71"),
   326 => (x"4f",x"26",x"58",x"f5"),
   327 => (x"5c",x"5b",x"5e",x"0e"),
   328 => (x"4b",x"71",x"0e",x"5d"),
   329 => (x"c2",x"87",x"c7",x"ff"),
   330 => (x"c0",x"48",x"e8",x"f6"),
   331 => (x"ff",x"49",x"73",x"50"),
   332 => (x"70",x"87",x"fe",x"db"),
   333 => (x"9c",x"c2",x"4c",x"49"),
   334 => (x"cb",x"49",x"ee",x"cb"),
   335 => (x"49",x"70",x"87",x"cf"),
   336 => (x"e8",x"f6",x"c2",x"4d"),
   337 => (x"c1",x"05",x"bf",x"97"),
   338 => (x"66",x"d0",x"87",x"e4"),
   339 => (x"f1",x"f6",x"c2",x"49"),
   340 => (x"d7",x"05",x"99",x"bf"),
   341 => (x"49",x"66",x"d4",x"87"),
   342 => (x"bf",x"e9",x"f6",x"c2"),
   343 => (x"87",x"cc",x"05",x"99"),
   344 => (x"db",x"ff",x"49",x"73"),
   345 => (x"98",x"70",x"87",x"cb"),
   346 => (x"87",x"c2",x"c1",x"02"),
   347 => (x"fd",x"fd",x"4c",x"c1"),
   348 => (x"ca",x"49",x"75",x"87"),
   349 => (x"98",x"70",x"87",x"e3"),
   350 => (x"c2",x"87",x"c6",x"02"),
   351 => (x"c1",x"48",x"e8",x"f6"),
   352 => (x"e8",x"f6",x"c2",x"50"),
   353 => (x"c0",x"05",x"bf",x"97"),
   354 => (x"f6",x"c2",x"87",x"e4"),
   355 => (x"d0",x"49",x"bf",x"f1"),
   356 => (x"ff",x"05",x"99",x"66"),
   357 => (x"f6",x"c2",x"87",x"d6"),
   358 => (x"d4",x"49",x"bf",x"e9"),
   359 => (x"ff",x"05",x"99",x"66"),
   360 => (x"49",x"73",x"87",x"ca"),
   361 => (x"87",x"c9",x"da",x"ff"),
   362 => (x"fe",x"05",x"98",x"70"),
   363 => (x"48",x"74",x"87",x"fe"),
   364 => (x"0e",x"87",x"d7",x"fb"),
   365 => (x"5d",x"5c",x"5b",x"5e"),
   366 => (x"c0",x"86",x"f4",x"0e"),
   367 => (x"bf",x"ec",x"4c",x"4d"),
   368 => (x"48",x"a6",x"c4",x"7e"),
   369 => (x"bf",x"f5",x"f6",x"c2"),
   370 => (x"c0",x"1e",x"c1",x"78"),
   371 => (x"fd",x"49",x"c7",x"1e"),
   372 => (x"86",x"c8",x"87",x"ca"),
   373 => (x"ce",x"02",x"98",x"70"),
   374 => (x"fb",x"49",x"ff",x"87"),
   375 => (x"da",x"c1",x"87",x"c7"),
   376 => (x"cc",x"d9",x"ff",x"49"),
   377 => (x"c2",x"4d",x"c1",x"87"),
   378 => (x"bf",x"97",x"e8",x"f6"),
   379 => (x"c9",x"87",x"c3",x"02"),
   380 => (x"f6",x"c2",x"87",x"c0"),
   381 => (x"c2",x"4b",x"bf",x"ed"),
   382 => (x"05",x"bf",x"c5",x"e0"),
   383 => (x"c3",x"87",x"eb",x"c0"),
   384 => (x"d8",x"ff",x"49",x"fd"),
   385 => (x"fa",x"c3",x"87",x"eb"),
   386 => (x"e4",x"d8",x"ff",x"49"),
   387 => (x"c3",x"49",x"73",x"87"),
   388 => (x"1e",x"71",x"99",x"ff"),
   389 => (x"c6",x"fb",x"49",x"c0"),
   390 => (x"c8",x"49",x"73",x"87"),
   391 => (x"1e",x"71",x"29",x"b7"),
   392 => (x"fa",x"fa",x"49",x"c1"),
   393 => (x"c6",x"86",x"c8",x"87"),
   394 => (x"f6",x"c2",x"87",x"c1"),
   395 => (x"9b",x"4b",x"bf",x"f1"),
   396 => (x"c2",x"87",x"dd",x"02"),
   397 => (x"49",x"bf",x"c1",x"e0"),
   398 => (x"70",x"87",x"de",x"c7"),
   399 => (x"87",x"c4",x"05",x"98"),
   400 => (x"87",x"d2",x"4b",x"c0"),
   401 => (x"c7",x"49",x"e0",x"c2"),
   402 => (x"e0",x"c2",x"87",x"c3"),
   403 => (x"87",x"c6",x"58",x"c5"),
   404 => (x"48",x"c1",x"e0",x"c2"),
   405 => (x"49",x"73",x"78",x"c0"),
   406 => (x"ce",x"05",x"99",x"c2"),
   407 => (x"49",x"eb",x"c3",x"87"),
   408 => (x"87",x"cd",x"d7",x"ff"),
   409 => (x"99",x"c2",x"49",x"70"),
   410 => (x"fb",x"87",x"c2",x"02"),
   411 => (x"c1",x"49",x"73",x"4c"),
   412 => (x"87",x"ce",x"05",x"99"),
   413 => (x"ff",x"49",x"f4",x"c3"),
   414 => (x"70",x"87",x"f6",x"d6"),
   415 => (x"02",x"99",x"c2",x"49"),
   416 => (x"4c",x"fa",x"87",x"c2"),
   417 => (x"99",x"c8",x"49",x"73"),
   418 => (x"c3",x"87",x"ce",x"05"),
   419 => (x"d6",x"ff",x"49",x"f5"),
   420 => (x"49",x"70",x"87",x"df"),
   421 => (x"d5",x"02",x"99",x"c2"),
   422 => (x"f9",x"f6",x"c2",x"87"),
   423 => (x"87",x"ca",x"02",x"bf"),
   424 => (x"c2",x"88",x"c1",x"48"),
   425 => (x"c0",x"58",x"fd",x"f6"),
   426 => (x"4c",x"ff",x"87",x"c2"),
   427 => (x"49",x"73",x"4d",x"c1"),
   428 => (x"ce",x"05",x"99",x"c4"),
   429 => (x"49",x"f2",x"c3",x"87"),
   430 => (x"87",x"f5",x"d5",x"ff"),
   431 => (x"99",x"c2",x"49",x"70"),
   432 => (x"c2",x"87",x"dc",x"02"),
   433 => (x"7e",x"bf",x"f9",x"f6"),
   434 => (x"a8",x"b7",x"c7",x"48"),
   435 => (x"87",x"cb",x"c0",x"03"),
   436 => (x"80",x"c1",x"48",x"6e"),
   437 => (x"58",x"fd",x"f6",x"c2"),
   438 => (x"fe",x"87",x"c2",x"c0"),
   439 => (x"c3",x"4d",x"c1",x"4c"),
   440 => (x"d5",x"ff",x"49",x"fd"),
   441 => (x"49",x"70",x"87",x"cb"),
   442 => (x"c0",x"02",x"99",x"c2"),
   443 => (x"f6",x"c2",x"87",x"d5"),
   444 => (x"c0",x"02",x"bf",x"f9"),
   445 => (x"f6",x"c2",x"87",x"c9"),
   446 => (x"78",x"c0",x"48",x"f9"),
   447 => (x"fd",x"87",x"c2",x"c0"),
   448 => (x"c3",x"4d",x"c1",x"4c"),
   449 => (x"d4",x"ff",x"49",x"fa"),
   450 => (x"49",x"70",x"87",x"e7"),
   451 => (x"c0",x"02",x"99",x"c2"),
   452 => (x"f6",x"c2",x"87",x"d9"),
   453 => (x"c7",x"48",x"bf",x"f9"),
   454 => (x"c0",x"03",x"a8",x"b7"),
   455 => (x"f6",x"c2",x"87",x"c9"),
   456 => (x"78",x"c7",x"48",x"f9"),
   457 => (x"fc",x"87",x"c2",x"c0"),
   458 => (x"c0",x"4d",x"c1",x"4c"),
   459 => (x"c0",x"03",x"ac",x"b7"),
   460 => (x"66",x"c4",x"87",x"d1"),
   461 => (x"82",x"d8",x"c1",x"4a"),
   462 => (x"c6",x"c0",x"02",x"6a"),
   463 => (x"74",x"4b",x"6a",x"87"),
   464 => (x"c0",x"0f",x"73",x"49"),
   465 => (x"1e",x"f0",x"c3",x"1e"),
   466 => (x"f7",x"49",x"da",x"c1"),
   467 => (x"86",x"c8",x"87",x"ce"),
   468 => (x"c0",x"02",x"98",x"70"),
   469 => (x"a6",x"c8",x"87",x"e2"),
   470 => (x"f9",x"f6",x"c2",x"48"),
   471 => (x"66",x"c8",x"78",x"bf"),
   472 => (x"c4",x"91",x"cb",x"49"),
   473 => (x"80",x"71",x"48",x"66"),
   474 => (x"bf",x"6e",x"7e",x"70"),
   475 => (x"87",x"c8",x"c0",x"02"),
   476 => (x"c8",x"4b",x"bf",x"6e"),
   477 => (x"0f",x"73",x"49",x"66"),
   478 => (x"c0",x"02",x"9d",x"75"),
   479 => (x"f6",x"c2",x"87",x"c8"),
   480 => (x"f2",x"49",x"bf",x"f9"),
   481 => (x"e0",x"c2",x"87",x"fa"),
   482 => (x"c0",x"02",x"bf",x"c9"),
   483 => (x"c2",x"49",x"87",x"dd"),
   484 => (x"98",x"70",x"87",x"c7"),
   485 => (x"87",x"d3",x"c0",x"02"),
   486 => (x"bf",x"f9",x"f6",x"c2"),
   487 => (x"87",x"e0",x"f2",x"49"),
   488 => (x"c0",x"f4",x"49",x"c0"),
   489 => (x"c9",x"e0",x"c2",x"87"),
   490 => (x"f4",x"78",x"c0",x"48"),
   491 => (x"87",x"da",x"f3",x"8e"),
   492 => (x"5c",x"5b",x"5e",x"0e"),
   493 => (x"71",x"1e",x"0e",x"5d"),
   494 => (x"f5",x"f6",x"c2",x"4c"),
   495 => (x"cd",x"c1",x"49",x"bf"),
   496 => (x"d1",x"c1",x"4d",x"a1"),
   497 => (x"74",x"7e",x"69",x"81"),
   498 => (x"87",x"cf",x"02",x"9c"),
   499 => (x"74",x"4b",x"a5",x"c4"),
   500 => (x"f5",x"f6",x"c2",x"7b"),
   501 => (x"f9",x"f2",x"49",x"bf"),
   502 => (x"74",x"7b",x"6e",x"87"),
   503 => (x"87",x"c4",x"05",x"9c"),
   504 => (x"87",x"c2",x"4b",x"c0"),
   505 => (x"49",x"73",x"4b",x"c1"),
   506 => (x"d4",x"87",x"fa",x"f2"),
   507 => (x"87",x"c7",x"02",x"66"),
   508 => (x"70",x"87",x"da",x"49"),
   509 => (x"c0",x"87",x"c2",x"4a"),
   510 => (x"cd",x"e0",x"c2",x"4a"),
   511 => (x"c9",x"f2",x"26",x"5a"),
   512 => (x"00",x"00",x"00",x"87"),
   513 => (x"00",x"00",x"00",x"00"),
   514 => (x"00",x"00",x"00",x"00"),
   515 => (x"4a",x"71",x"1e",x"00"),
   516 => (x"49",x"bf",x"c8",x"ff"),
   517 => (x"26",x"48",x"a1",x"72"),
   518 => (x"c8",x"ff",x"1e",x"4f"),
   519 => (x"c0",x"fe",x"89",x"bf"),
   520 => (x"c0",x"c0",x"c0",x"c0"),
   521 => (x"87",x"c4",x"01",x"a9"),
   522 => (x"87",x"c2",x"4a",x"c0"),
   523 => (x"48",x"72",x"4a",x"c1"),
   524 => (x"c2",x"1e",x"4f",x"26"),
   525 => (x"49",x"bf",x"db",x"e1"),
   526 => (x"e1",x"c2",x"b9",x"c1"),
   527 => (x"d4",x"ff",x"59",x"df"),
   528 => (x"78",x"ff",x"c3",x"48"),
   529 => (x"c0",x"48",x"d0",x"ff"),
   530 => (x"d4",x"ff",x"78",x"e1"),
   531 => (x"c4",x"78",x"c1",x"48"),
   532 => (x"ff",x"78",x"71",x"31"),
   533 => (x"e0",x"c0",x"48",x"d0"),
   534 => (x"00",x"4f",x"26",x"78"),
   535 => (x"0e",x"00",x"00",x"00"),
   536 => (x"5d",x"5c",x"5b",x"5e"),
   537 => (x"e9",x"f6",x"c2",x"0e"),
   538 => (x"e3",x"c2",x"4a",x"bf"),
   539 => (x"4c",x"49",x"bf",x"c8"),
   540 => (x"4d",x"71",x"bc",x"72"),
   541 => (x"87",x"e0",x"c7",x"ff"),
   542 => (x"49",x"74",x"4b",x"c0"),
   543 => (x"c0",x"02",x"99",x"d0"),
   544 => (x"d0",x"ff",x"87",x"e7"),
   545 => (x"78",x"e1",x"c8",x"48"),
   546 => (x"c5",x"48",x"d4",x"ff"),
   547 => (x"d0",x"49",x"75",x"78"),
   548 => (x"87",x"c3",x"02",x"99"),
   549 => (x"c2",x"78",x"f0",x"c3"),
   550 => (x"73",x"49",x"f6",x"e3"),
   551 => (x"ff",x"48",x"11",x"81"),
   552 => (x"ff",x"78",x"08",x"d4"),
   553 => (x"e0",x"c0",x"48",x"d0"),
   554 => (x"2d",x"2c",x"c1",x"78"),
   555 => (x"04",x"ab",x"c8",x"83"),
   556 => (x"ff",x"87",x"c7",x"ff"),
   557 => (x"c2",x"87",x"d9",x"c6"),
   558 => (x"c2",x"48",x"c8",x"e3"),
   559 => (x"78",x"bf",x"e9",x"f6"),
   560 => (x"4c",x"26",x"4d",x"26"),
   561 => (x"4f",x"26",x"4b",x"26"),
   562 => (x"00",x"00",x"00",x"00"),
   563 => (x"c3",x"e7",x"c1",x"1e"),
   564 => (x"c2",x"50",x"de",x"48"),
   565 => (x"fe",x"49",x"df",x"e3"),
   566 => (x"c0",x"87",x"ea",x"da"),
   567 => (x"50",x"4f",x"26",x"48"),
   568 => (x"4d",x"4b",x"43",x"55"),
   569 => (x"41",x"31",x"7e",x"41"),
   570 => (x"1e",x"00",x"43",x"52"),
   571 => (x"fd",x"87",x"c4",x"f3"),
   572 => (x"87",x"f8",x"87",x"ed"),
   573 => (x"1e",x"16",x"4f",x"26"),
   574 => (x"36",x"2e",x"25",x"26"),
   575 => (x"36",x"2e",x"3e",x"3d"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

