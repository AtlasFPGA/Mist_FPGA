
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"c0",x"f7",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"c0",x"f7",x"c2"),
    14 => (x"48",x"c0",x"e4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"e0",x"e5"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"81",x"48",x"73",x"1e"),
    47 => (x"72",x"05",x"a9",x"73"),
    48 => (x"26",x"87",x"f9",x"53"),
    49 => (x"4a",x"71",x"1e",x"4f"),
    50 => (x"48",x"49",x"66",x"c4"),
    51 => (x"a6",x"c8",x"88",x"c1"),
    52 => (x"02",x"99",x"71",x"58"),
    53 => (x"d4",x"ff",x"87",x"d6"),
    54 => (x"78",x"ff",x"c3",x"48"),
    55 => (x"66",x"c4",x"52",x"68"),
    56 => (x"88",x"c1",x"48",x"49"),
    57 => (x"71",x"58",x"a6",x"c8"),
    58 => (x"87",x"ea",x"05",x"99"),
    59 => (x"73",x"1e",x"4f",x"26"),
    60 => (x"4b",x"d4",x"ff",x"1e"),
    61 => (x"6b",x"7b",x"ff",x"c3"),
    62 => (x"7b",x"ff",x"c3",x"4a"),
    63 => (x"32",x"c8",x"49",x"6b"),
    64 => (x"ff",x"c3",x"b1",x"72"),
    65 => (x"c8",x"4a",x"6b",x"7b"),
    66 => (x"c3",x"b2",x"71",x"31"),
    67 => (x"49",x"6b",x"7b",x"ff"),
    68 => (x"b1",x"72",x"32",x"c8"),
    69 => (x"87",x"c4",x"48",x"71"),
    70 => (x"4c",x"26",x"4d",x"26"),
    71 => (x"4f",x"26",x"4b",x"26"),
    72 => (x"5c",x"5b",x"5e",x"0e"),
    73 => (x"4a",x"71",x"0e",x"5d"),
    74 => (x"72",x"4c",x"d4",x"ff"),
    75 => (x"99",x"ff",x"c3",x"49"),
    76 => (x"e4",x"c2",x"7c",x"71"),
    77 => (x"c8",x"05",x"bf",x"c0"),
    78 => (x"48",x"66",x"d0",x"87"),
    79 => (x"a6",x"d4",x"30",x"c9"),
    80 => (x"49",x"66",x"d0",x"58"),
    81 => (x"ff",x"c3",x"29",x"d8"),
    82 => (x"d0",x"7c",x"71",x"99"),
    83 => (x"29",x"d0",x"49",x"66"),
    84 => (x"71",x"99",x"ff",x"c3"),
    85 => (x"49",x"66",x"d0",x"7c"),
    86 => (x"ff",x"c3",x"29",x"c8"),
    87 => (x"d0",x"7c",x"71",x"99"),
    88 => (x"ff",x"c3",x"49",x"66"),
    89 => (x"72",x"7c",x"71",x"99"),
    90 => (x"c3",x"29",x"d0",x"49"),
    91 => (x"7c",x"71",x"99",x"ff"),
    92 => (x"f0",x"c9",x"4b",x"6c"),
    93 => (x"ff",x"c3",x"4d",x"ff"),
    94 => (x"87",x"d0",x"05",x"ab"),
    95 => (x"6c",x"7c",x"ff",x"c3"),
    96 => (x"02",x"8d",x"c1",x"4b"),
    97 => (x"ff",x"c3",x"87",x"c6"),
    98 => (x"87",x"f0",x"02",x"ab"),
    99 => (x"c7",x"fe",x"48",x"73"),
   100 => (x"49",x"c0",x"1e",x"87"),
   101 => (x"c3",x"48",x"d4",x"ff"),
   102 => (x"81",x"c1",x"78",x"ff"),
   103 => (x"a9",x"b7",x"c8",x"c3"),
   104 => (x"26",x"87",x"f1",x"04"),
   105 => (x"1e",x"73",x"1e",x"4f"),
   106 => (x"f8",x"c4",x"87",x"e7"),
   107 => (x"1e",x"c0",x"4b",x"df"),
   108 => (x"c1",x"f0",x"ff",x"c0"),
   109 => (x"e7",x"fd",x"49",x"f7"),
   110 => (x"c1",x"86",x"c4",x"87"),
   111 => (x"ea",x"c0",x"05",x"a8"),
   112 => (x"48",x"d4",x"ff",x"87"),
   113 => (x"c1",x"78",x"ff",x"c3"),
   114 => (x"c0",x"c0",x"c0",x"c0"),
   115 => (x"e1",x"c0",x"1e",x"c0"),
   116 => (x"49",x"e9",x"c1",x"f0"),
   117 => (x"c4",x"87",x"c9",x"fd"),
   118 => (x"05",x"98",x"70",x"86"),
   119 => (x"d4",x"ff",x"87",x"ca"),
   120 => (x"78",x"ff",x"c3",x"48"),
   121 => (x"87",x"cb",x"48",x"c1"),
   122 => (x"c1",x"87",x"e6",x"fe"),
   123 => (x"fd",x"fe",x"05",x"8b"),
   124 => (x"fc",x"48",x"c0",x"87"),
   125 => (x"73",x"1e",x"87",x"e6"),
   126 => (x"48",x"d4",x"ff",x"1e"),
   127 => (x"d3",x"78",x"ff",x"c3"),
   128 => (x"c0",x"1e",x"c0",x"4b"),
   129 => (x"c1",x"c1",x"f0",x"ff"),
   130 => (x"87",x"d4",x"fc",x"49"),
   131 => (x"98",x"70",x"86",x"c4"),
   132 => (x"ff",x"87",x"ca",x"05"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"cb",x"48",x"c1",x"78"),
   135 => (x"87",x"f1",x"fd",x"87"),
   136 => (x"ff",x"05",x"8b",x"c1"),
   137 => (x"48",x"c0",x"87",x"db"),
   138 => (x"0e",x"87",x"f1",x"fb"),
   139 => (x"0e",x"5c",x"5b",x"5e"),
   140 => (x"fd",x"4c",x"d4",x"ff"),
   141 => (x"ea",x"c6",x"87",x"db"),
   142 => (x"f0",x"e1",x"c0",x"1e"),
   143 => (x"fb",x"49",x"c8",x"c1"),
   144 => (x"86",x"c4",x"87",x"de"),
   145 => (x"c8",x"02",x"a8",x"c1"),
   146 => (x"87",x"ea",x"fe",x"87"),
   147 => (x"e2",x"c1",x"48",x"c0"),
   148 => (x"87",x"da",x"fa",x"87"),
   149 => (x"ff",x"cf",x"49",x"70"),
   150 => (x"ea",x"c6",x"99",x"ff"),
   151 => (x"87",x"c8",x"02",x"a9"),
   152 => (x"c0",x"87",x"d3",x"fe"),
   153 => (x"87",x"cb",x"c1",x"48"),
   154 => (x"c0",x"7c",x"ff",x"c3"),
   155 => (x"f4",x"fc",x"4b",x"f1"),
   156 => (x"02",x"98",x"70",x"87"),
   157 => (x"c0",x"87",x"eb",x"c0"),
   158 => (x"f0",x"ff",x"c0",x"1e"),
   159 => (x"fa",x"49",x"fa",x"c1"),
   160 => (x"86",x"c4",x"87",x"de"),
   161 => (x"d9",x"05",x"98",x"70"),
   162 => (x"7c",x"ff",x"c3",x"87"),
   163 => (x"ff",x"c3",x"49",x"6c"),
   164 => (x"7c",x"7c",x"7c",x"7c"),
   165 => (x"02",x"99",x"c0",x"c1"),
   166 => (x"48",x"c1",x"87",x"c4"),
   167 => (x"48",x"c0",x"87",x"d5"),
   168 => (x"ab",x"c2",x"87",x"d1"),
   169 => (x"c0",x"87",x"c4",x"05"),
   170 => (x"c1",x"87",x"c8",x"48"),
   171 => (x"fd",x"fe",x"05",x"8b"),
   172 => (x"f9",x"48",x"c0",x"87"),
   173 => (x"73",x"1e",x"87",x"e4"),
   174 => (x"c0",x"e4",x"c2",x"1e"),
   175 => (x"c7",x"78",x"c1",x"48"),
   176 => (x"48",x"d0",x"ff",x"4b"),
   177 => (x"c8",x"fb",x"78",x"c2"),
   178 => (x"48",x"d0",x"ff",x"87"),
   179 => (x"1e",x"c0",x"78",x"c3"),
   180 => (x"c1",x"d0",x"e5",x"c0"),
   181 => (x"c7",x"f9",x"49",x"c0"),
   182 => (x"c1",x"86",x"c4",x"87"),
   183 => (x"87",x"c1",x"05",x"a8"),
   184 => (x"05",x"ab",x"c2",x"4b"),
   185 => (x"48",x"c0",x"87",x"c5"),
   186 => (x"c1",x"87",x"f9",x"c0"),
   187 => (x"d0",x"ff",x"05",x"8b"),
   188 => (x"87",x"f7",x"fc",x"87"),
   189 => (x"58",x"c4",x"e4",x"c2"),
   190 => (x"cd",x"05",x"98",x"70"),
   191 => (x"c0",x"1e",x"c1",x"87"),
   192 => (x"d0",x"c1",x"f0",x"ff"),
   193 => (x"87",x"d8",x"f8",x"49"),
   194 => (x"d4",x"ff",x"86",x"c4"),
   195 => (x"78",x"ff",x"c3",x"48"),
   196 => (x"c2",x"87",x"fc",x"c2"),
   197 => (x"ff",x"58",x"c8",x"e4"),
   198 => (x"78",x"c2",x"48",x"d0"),
   199 => (x"c3",x"48",x"d4",x"ff"),
   200 => (x"48",x"c1",x"78",x"ff"),
   201 => (x"0e",x"87",x"f5",x"f7"),
   202 => (x"5d",x"5c",x"5b",x"5e"),
   203 => (x"c0",x"4b",x"71",x"0e"),
   204 => (x"cd",x"ee",x"c5",x"4c"),
   205 => (x"d4",x"ff",x"4a",x"df"),
   206 => (x"78",x"ff",x"c3",x"48"),
   207 => (x"fe",x"c3",x"49",x"68"),
   208 => (x"fd",x"c0",x"05",x"a9"),
   209 => (x"73",x"4d",x"70",x"87"),
   210 => (x"87",x"cc",x"02",x"9b"),
   211 => (x"73",x"1e",x"66",x"d0"),
   212 => (x"87",x"f1",x"f5",x"49"),
   213 => (x"87",x"d6",x"86",x"c4"),
   214 => (x"c4",x"48",x"d0",x"ff"),
   215 => (x"ff",x"c3",x"78",x"d1"),
   216 => (x"48",x"66",x"d0",x"7d"),
   217 => (x"a6",x"d4",x"88",x"c1"),
   218 => (x"05",x"98",x"70",x"58"),
   219 => (x"d4",x"ff",x"87",x"f0"),
   220 => (x"78",x"ff",x"c3",x"48"),
   221 => (x"05",x"9b",x"73",x"78"),
   222 => (x"d0",x"ff",x"87",x"c5"),
   223 => (x"c1",x"78",x"d0",x"48"),
   224 => (x"8a",x"c1",x"4c",x"4a"),
   225 => (x"87",x"ee",x"fe",x"05"),
   226 => (x"cb",x"f6",x"48",x"74"),
   227 => (x"1e",x"73",x"1e",x"87"),
   228 => (x"4b",x"c0",x"4a",x"71"),
   229 => (x"c3",x"48",x"d4",x"ff"),
   230 => (x"d0",x"ff",x"78",x"ff"),
   231 => (x"78",x"c3",x"c4",x"48"),
   232 => (x"c3",x"48",x"d4",x"ff"),
   233 => (x"1e",x"72",x"78",x"ff"),
   234 => (x"c1",x"f0",x"ff",x"c0"),
   235 => (x"ef",x"f5",x"49",x"d1"),
   236 => (x"70",x"86",x"c4",x"87"),
   237 => (x"87",x"d2",x"05",x"98"),
   238 => (x"cc",x"1e",x"c0",x"c8"),
   239 => (x"e6",x"fd",x"49",x"66"),
   240 => (x"70",x"86",x"c4",x"87"),
   241 => (x"48",x"d0",x"ff",x"4b"),
   242 => (x"48",x"73",x"78",x"c2"),
   243 => (x"0e",x"87",x"cd",x"f5"),
   244 => (x"5d",x"5c",x"5b",x"5e"),
   245 => (x"c0",x"1e",x"c0",x"0e"),
   246 => (x"c9",x"c1",x"f0",x"ff"),
   247 => (x"87",x"c0",x"f5",x"49"),
   248 => (x"e4",x"c2",x"1e",x"d2"),
   249 => (x"fe",x"fc",x"49",x"c8"),
   250 => (x"c0",x"86",x"c8",x"87"),
   251 => (x"d2",x"84",x"c1",x"4c"),
   252 => (x"f8",x"04",x"ac",x"b7"),
   253 => (x"c8",x"e4",x"c2",x"87"),
   254 => (x"c3",x"49",x"bf",x"97"),
   255 => (x"c0",x"c1",x"99",x"c0"),
   256 => (x"e7",x"c0",x"05",x"a9"),
   257 => (x"cf",x"e4",x"c2",x"87"),
   258 => (x"d0",x"49",x"bf",x"97"),
   259 => (x"d0",x"e4",x"c2",x"31"),
   260 => (x"c8",x"4a",x"bf",x"97"),
   261 => (x"c2",x"b1",x"72",x"32"),
   262 => (x"bf",x"97",x"d1",x"e4"),
   263 => (x"4c",x"71",x"b1",x"4a"),
   264 => (x"ff",x"ff",x"ff",x"cf"),
   265 => (x"ca",x"84",x"c1",x"9c"),
   266 => (x"87",x"e7",x"c1",x"34"),
   267 => (x"97",x"d1",x"e4",x"c2"),
   268 => (x"31",x"c1",x"49",x"bf"),
   269 => (x"e4",x"c2",x"99",x"c6"),
   270 => (x"4a",x"bf",x"97",x"d2"),
   271 => (x"72",x"2a",x"b7",x"c7"),
   272 => (x"cd",x"e4",x"c2",x"b1"),
   273 => (x"4d",x"4a",x"bf",x"97"),
   274 => (x"e4",x"c2",x"9d",x"cf"),
   275 => (x"4a",x"bf",x"97",x"ce"),
   276 => (x"32",x"ca",x"9a",x"c3"),
   277 => (x"97",x"cf",x"e4",x"c2"),
   278 => (x"33",x"c2",x"4b",x"bf"),
   279 => (x"e4",x"c2",x"b2",x"73"),
   280 => (x"4b",x"bf",x"97",x"d0"),
   281 => (x"c6",x"9b",x"c0",x"c3"),
   282 => (x"b2",x"73",x"2b",x"b7"),
   283 => (x"48",x"c1",x"81",x"c2"),
   284 => (x"49",x"70",x"30",x"71"),
   285 => (x"30",x"75",x"48",x"c1"),
   286 => (x"4c",x"72",x"4d",x"70"),
   287 => (x"94",x"71",x"84",x"c1"),
   288 => (x"ad",x"b7",x"c0",x"c8"),
   289 => (x"c1",x"87",x"cc",x"06"),
   290 => (x"c8",x"2d",x"b7",x"34"),
   291 => (x"01",x"ad",x"b7",x"c0"),
   292 => (x"74",x"87",x"f4",x"ff"),
   293 => (x"87",x"c0",x"f2",x"48"),
   294 => (x"5c",x"5b",x"5e",x"0e"),
   295 => (x"86",x"f8",x"0e",x"5d"),
   296 => (x"48",x"ee",x"ec",x"c2"),
   297 => (x"e4",x"c2",x"78",x"c0"),
   298 => (x"49",x"c0",x"1e",x"e6"),
   299 => (x"c4",x"87",x"de",x"fb"),
   300 => (x"05",x"98",x"70",x"86"),
   301 => (x"48",x"c0",x"87",x"c5"),
   302 => (x"c0",x"87",x"ce",x"c9"),
   303 => (x"c0",x"7e",x"c1",x"4d"),
   304 => (x"49",x"bf",x"cf",x"f5"),
   305 => (x"4a",x"dc",x"e5",x"c2"),
   306 => (x"ee",x"4b",x"c8",x"71"),
   307 => (x"98",x"70",x"87",x"dc"),
   308 => (x"c0",x"87",x"c2",x"05"),
   309 => (x"cb",x"f5",x"c0",x"7e"),
   310 => (x"e5",x"c2",x"49",x"bf"),
   311 => (x"c8",x"71",x"4a",x"f8"),
   312 => (x"87",x"c6",x"ee",x"4b"),
   313 => (x"c2",x"05",x"98",x"70"),
   314 => (x"6e",x"7e",x"c0",x"87"),
   315 => (x"87",x"fd",x"c0",x"02"),
   316 => (x"bf",x"ec",x"eb",x"c2"),
   317 => (x"e4",x"ec",x"c2",x"4d"),
   318 => (x"48",x"7e",x"bf",x"9f"),
   319 => (x"a8",x"ea",x"d6",x"c5"),
   320 => (x"c2",x"87",x"c7",x"05"),
   321 => (x"4d",x"bf",x"ec",x"eb"),
   322 => (x"48",x"6e",x"87",x"ce"),
   323 => (x"a8",x"d5",x"e9",x"ca"),
   324 => (x"c0",x"87",x"c5",x"02"),
   325 => (x"87",x"f1",x"c7",x"48"),
   326 => (x"1e",x"e6",x"e4",x"c2"),
   327 => (x"ec",x"f9",x"49",x"75"),
   328 => (x"70",x"86",x"c4",x"87"),
   329 => (x"87",x"c5",x"05",x"98"),
   330 => (x"dc",x"c7",x"48",x"c0"),
   331 => (x"cb",x"f5",x"c0",x"87"),
   332 => (x"e5",x"c2",x"49",x"bf"),
   333 => (x"c8",x"71",x"4a",x"f8"),
   334 => (x"87",x"ee",x"ec",x"4b"),
   335 => (x"c8",x"05",x"98",x"70"),
   336 => (x"ee",x"ec",x"c2",x"87"),
   337 => (x"da",x"78",x"c1",x"48"),
   338 => (x"cf",x"f5",x"c0",x"87"),
   339 => (x"e5",x"c2",x"49",x"bf"),
   340 => (x"c8",x"71",x"4a",x"dc"),
   341 => (x"87",x"d2",x"ec",x"4b"),
   342 => (x"c0",x"02",x"98",x"70"),
   343 => (x"48",x"c0",x"87",x"c5"),
   344 => (x"c2",x"87",x"e6",x"c6"),
   345 => (x"bf",x"97",x"e4",x"ec"),
   346 => (x"a9",x"d5",x"c1",x"49"),
   347 => (x"87",x"cd",x"c0",x"05"),
   348 => (x"97",x"e5",x"ec",x"c2"),
   349 => (x"ea",x"c2",x"49",x"bf"),
   350 => (x"c5",x"c0",x"02",x"a9"),
   351 => (x"c6",x"48",x"c0",x"87"),
   352 => (x"e4",x"c2",x"87",x"c7"),
   353 => (x"7e",x"bf",x"97",x"e6"),
   354 => (x"a8",x"e9",x"c3",x"48"),
   355 => (x"87",x"ce",x"c0",x"02"),
   356 => (x"eb",x"c3",x"48",x"6e"),
   357 => (x"c5",x"c0",x"02",x"a8"),
   358 => (x"c5",x"48",x"c0",x"87"),
   359 => (x"e4",x"c2",x"87",x"eb"),
   360 => (x"49",x"bf",x"97",x"f1"),
   361 => (x"cc",x"c0",x"05",x"99"),
   362 => (x"f2",x"e4",x"c2",x"87"),
   363 => (x"c2",x"49",x"bf",x"97"),
   364 => (x"c5",x"c0",x"02",x"a9"),
   365 => (x"c5",x"48",x"c0",x"87"),
   366 => (x"e4",x"c2",x"87",x"cf"),
   367 => (x"48",x"bf",x"97",x"f3"),
   368 => (x"58",x"ea",x"ec",x"c2"),
   369 => (x"c1",x"48",x"4c",x"70"),
   370 => (x"ee",x"ec",x"c2",x"88"),
   371 => (x"f4",x"e4",x"c2",x"58"),
   372 => (x"75",x"49",x"bf",x"97"),
   373 => (x"f5",x"e4",x"c2",x"81"),
   374 => (x"c8",x"4a",x"bf",x"97"),
   375 => (x"7e",x"a1",x"72",x"32"),
   376 => (x"48",x"fb",x"f0",x"c2"),
   377 => (x"e4",x"c2",x"78",x"6e"),
   378 => (x"48",x"bf",x"97",x"f6"),
   379 => (x"c2",x"58",x"a6",x"c8"),
   380 => (x"02",x"bf",x"ee",x"ec"),
   381 => (x"c0",x"87",x"d4",x"c2"),
   382 => (x"49",x"bf",x"cb",x"f5"),
   383 => (x"4a",x"f8",x"e5",x"c2"),
   384 => (x"e9",x"4b",x"c8",x"71"),
   385 => (x"98",x"70",x"87",x"e4"),
   386 => (x"87",x"c5",x"c0",x"02"),
   387 => (x"f8",x"c3",x"48",x"c0"),
   388 => (x"e6",x"ec",x"c2",x"87"),
   389 => (x"f1",x"c2",x"4c",x"bf"),
   390 => (x"e5",x"c2",x"5c",x"cf"),
   391 => (x"49",x"bf",x"97",x"cb"),
   392 => (x"e5",x"c2",x"31",x"c8"),
   393 => (x"4a",x"bf",x"97",x"ca"),
   394 => (x"e5",x"c2",x"49",x"a1"),
   395 => (x"4a",x"bf",x"97",x"cc"),
   396 => (x"a1",x"72",x"32",x"d0"),
   397 => (x"cd",x"e5",x"c2",x"49"),
   398 => (x"d8",x"4a",x"bf",x"97"),
   399 => (x"49",x"a1",x"72",x"32"),
   400 => (x"c2",x"91",x"66",x"c4"),
   401 => (x"81",x"bf",x"fb",x"f0"),
   402 => (x"59",x"c3",x"f1",x"c2"),
   403 => (x"97",x"d3",x"e5",x"c2"),
   404 => (x"32",x"c8",x"4a",x"bf"),
   405 => (x"97",x"d2",x"e5",x"c2"),
   406 => (x"4a",x"a2",x"4b",x"bf"),
   407 => (x"97",x"d4",x"e5",x"c2"),
   408 => (x"33",x"d0",x"4b",x"bf"),
   409 => (x"c2",x"4a",x"a2",x"73"),
   410 => (x"bf",x"97",x"d5",x"e5"),
   411 => (x"d8",x"9b",x"cf",x"4b"),
   412 => (x"4a",x"a2",x"73",x"33"),
   413 => (x"5a",x"c7",x"f1",x"c2"),
   414 => (x"bf",x"c3",x"f1",x"c2"),
   415 => (x"74",x"8a",x"c2",x"4a"),
   416 => (x"c7",x"f1",x"c2",x"92"),
   417 => (x"78",x"a1",x"72",x"48"),
   418 => (x"c2",x"87",x"ca",x"c1"),
   419 => (x"bf",x"97",x"f8",x"e4"),
   420 => (x"c2",x"31",x"c8",x"49"),
   421 => (x"bf",x"97",x"f7",x"e4"),
   422 => (x"c2",x"49",x"a1",x"4a"),
   423 => (x"c2",x"59",x"f6",x"ec"),
   424 => (x"49",x"bf",x"f2",x"ec"),
   425 => (x"ff",x"c7",x"31",x"c5"),
   426 => (x"c2",x"29",x"c9",x"81"),
   427 => (x"c2",x"59",x"cf",x"f1"),
   428 => (x"bf",x"97",x"fd",x"e4"),
   429 => (x"c2",x"32",x"c8",x"4a"),
   430 => (x"bf",x"97",x"fc",x"e4"),
   431 => (x"c4",x"4a",x"a2",x"4b"),
   432 => (x"82",x"6e",x"92",x"66"),
   433 => (x"5a",x"cb",x"f1",x"c2"),
   434 => (x"48",x"c3",x"f1",x"c2"),
   435 => (x"f0",x"c2",x"78",x"c0"),
   436 => (x"a1",x"72",x"48",x"ff"),
   437 => (x"cf",x"f1",x"c2",x"78"),
   438 => (x"c3",x"f1",x"c2",x"48"),
   439 => (x"f1",x"c2",x"78",x"bf"),
   440 => (x"f1",x"c2",x"48",x"d3"),
   441 => (x"c2",x"78",x"bf",x"c7"),
   442 => (x"02",x"bf",x"ee",x"ec"),
   443 => (x"74",x"87",x"c9",x"c0"),
   444 => (x"70",x"30",x"c4",x"48"),
   445 => (x"87",x"c9",x"c0",x"7e"),
   446 => (x"bf",x"cb",x"f1",x"c2"),
   447 => (x"70",x"30",x"c4",x"48"),
   448 => (x"f2",x"ec",x"c2",x"7e"),
   449 => (x"c1",x"78",x"6e",x"48"),
   450 => (x"26",x"8e",x"f8",x"48"),
   451 => (x"26",x"4c",x"26",x"4d"),
   452 => (x"0e",x"4f",x"26",x"4b"),
   453 => (x"5d",x"5c",x"5b",x"5e"),
   454 => (x"c2",x"4a",x"71",x"0e"),
   455 => (x"02",x"bf",x"ee",x"ec"),
   456 => (x"4b",x"72",x"87",x"cb"),
   457 => (x"4c",x"72",x"2b",x"c7"),
   458 => (x"c9",x"9c",x"ff",x"c1"),
   459 => (x"c8",x"4b",x"72",x"87"),
   460 => (x"c3",x"4c",x"72",x"2b"),
   461 => (x"f0",x"c2",x"9c",x"ff"),
   462 => (x"c0",x"83",x"bf",x"fb"),
   463 => (x"ab",x"bf",x"c7",x"f5"),
   464 => (x"c0",x"87",x"d9",x"02"),
   465 => (x"c2",x"5b",x"cb",x"f5"),
   466 => (x"73",x"1e",x"e6",x"e4"),
   467 => (x"87",x"fd",x"f0",x"49"),
   468 => (x"98",x"70",x"86",x"c4"),
   469 => (x"c0",x"87",x"c5",x"05"),
   470 => (x"87",x"e6",x"c0",x"48"),
   471 => (x"bf",x"ee",x"ec",x"c2"),
   472 => (x"74",x"87",x"d2",x"02"),
   473 => (x"c2",x"91",x"c4",x"49"),
   474 => (x"69",x"81",x"e6",x"e4"),
   475 => (x"ff",x"ff",x"cf",x"4d"),
   476 => (x"cb",x"9d",x"ff",x"ff"),
   477 => (x"c2",x"49",x"74",x"87"),
   478 => (x"e6",x"e4",x"c2",x"91"),
   479 => (x"4d",x"69",x"9f",x"81"),
   480 => (x"c6",x"fe",x"48",x"75"),
   481 => (x"5b",x"5e",x"0e",x"87"),
   482 => (x"f8",x"0e",x"5d",x"5c"),
   483 => (x"9c",x"4c",x"71",x"86"),
   484 => (x"c0",x"87",x"c5",x"05"),
   485 => (x"87",x"c1",x"c3",x"48"),
   486 => (x"6e",x"7e",x"a4",x"c8"),
   487 => (x"d8",x"78",x"c0",x"48"),
   488 => (x"87",x"c7",x"02",x"66"),
   489 => (x"bf",x"97",x"66",x"d8"),
   490 => (x"c0",x"87",x"c5",x"05"),
   491 => (x"87",x"e9",x"c2",x"48"),
   492 => (x"49",x"c1",x"1e",x"c0"),
   493 => (x"c4",x"87",x"f4",x"ce"),
   494 => (x"9d",x"4d",x"70",x"86"),
   495 => (x"87",x"c2",x"c1",x"02"),
   496 => (x"4a",x"f6",x"ec",x"c2"),
   497 => (x"e2",x"49",x"66",x"d8"),
   498 => (x"98",x"70",x"87",x"c5"),
   499 => (x"87",x"f2",x"c0",x"02"),
   500 => (x"66",x"d8",x"4a",x"75"),
   501 => (x"e2",x"4b",x"cb",x"49"),
   502 => (x"98",x"70",x"87",x"ea"),
   503 => (x"87",x"e2",x"c0",x"02"),
   504 => (x"9d",x"75",x"1e",x"c0"),
   505 => (x"c8",x"87",x"c7",x"02"),
   506 => (x"78",x"c0",x"48",x"a6"),
   507 => (x"a6",x"c8",x"87",x"c5"),
   508 => (x"c8",x"78",x"c1",x"48"),
   509 => (x"f2",x"cd",x"49",x"66"),
   510 => (x"70",x"86",x"c4",x"87"),
   511 => (x"fe",x"05",x"9d",x"4d"),
   512 => (x"9d",x"75",x"87",x"fe"),
   513 => (x"87",x"cf",x"c1",x"02"),
   514 => (x"6e",x"49",x"a5",x"dc"),
   515 => (x"da",x"78",x"69",x"48"),
   516 => (x"a6",x"c4",x"49",x"a5"),
   517 => (x"78",x"a4",x"c4",x"48"),
   518 => (x"c4",x"48",x"69",x"9f"),
   519 => (x"c2",x"78",x"08",x"66"),
   520 => (x"02",x"bf",x"ee",x"ec"),
   521 => (x"a5",x"d4",x"87",x"d2"),
   522 => (x"49",x"69",x"9f",x"49"),
   523 => (x"99",x"ff",x"ff",x"c0"),
   524 => (x"30",x"d0",x"48",x"71"),
   525 => (x"87",x"c2",x"7e",x"70"),
   526 => (x"49",x"6e",x"7e",x"c0"),
   527 => (x"bf",x"66",x"c4",x"48"),
   528 => (x"08",x"66",x"c4",x"80"),
   529 => (x"cc",x"7c",x"c0",x"78"),
   530 => (x"66",x"c4",x"49",x"a4"),
   531 => (x"a4",x"d0",x"79",x"bf"),
   532 => (x"c1",x"79",x"c0",x"49"),
   533 => (x"c0",x"87",x"c2",x"48"),
   534 => (x"fa",x"8e",x"f8",x"48"),
   535 => (x"5e",x"0e",x"87",x"ed"),
   536 => (x"0e",x"5d",x"5c",x"5b"),
   537 => (x"02",x"9c",x"4c",x"71"),
   538 => (x"c8",x"87",x"ca",x"c1"),
   539 => (x"02",x"69",x"49",x"a4"),
   540 => (x"d0",x"87",x"c2",x"c1"),
   541 => (x"49",x"6c",x"4a",x"66"),
   542 => (x"5a",x"a6",x"d4",x"82"),
   543 => (x"b9",x"4d",x"66",x"d0"),
   544 => (x"bf",x"ea",x"ec",x"c2"),
   545 => (x"72",x"ba",x"ff",x"4a"),
   546 => (x"02",x"99",x"71",x"99"),
   547 => (x"c4",x"87",x"e4",x"c0"),
   548 => (x"49",x"6b",x"4b",x"a4"),
   549 => (x"70",x"87",x"fc",x"f9"),
   550 => (x"e6",x"ec",x"c2",x"7b"),
   551 => (x"81",x"6c",x"49",x"bf"),
   552 => (x"b9",x"75",x"7c",x"71"),
   553 => (x"bf",x"ea",x"ec",x"c2"),
   554 => (x"72",x"ba",x"ff",x"4a"),
   555 => (x"05",x"99",x"71",x"99"),
   556 => (x"75",x"87",x"dc",x"ff"),
   557 => (x"87",x"d3",x"f9",x"7c"),
   558 => (x"71",x"1e",x"73",x"1e"),
   559 => (x"c7",x"02",x"9b",x"4b"),
   560 => (x"49",x"a3",x"c8",x"87"),
   561 => (x"87",x"c5",x"05",x"69"),
   562 => (x"f7",x"c0",x"48",x"c0"),
   563 => (x"ff",x"f0",x"c2",x"87"),
   564 => (x"a3",x"c4",x"4a",x"bf"),
   565 => (x"c2",x"49",x"69",x"49"),
   566 => (x"e6",x"ec",x"c2",x"89"),
   567 => (x"a2",x"71",x"91",x"bf"),
   568 => (x"ea",x"ec",x"c2",x"4a"),
   569 => (x"99",x"6b",x"49",x"bf"),
   570 => (x"c0",x"4a",x"a2",x"71"),
   571 => (x"c8",x"5a",x"cb",x"f5"),
   572 => (x"49",x"72",x"1e",x"66"),
   573 => (x"c4",x"87",x"d6",x"ea"),
   574 => (x"05",x"98",x"70",x"86"),
   575 => (x"48",x"c0",x"87",x"c4"),
   576 => (x"48",x"c1",x"87",x"c2"),
   577 => (x"0e",x"87",x"c8",x"f8"),
   578 => (x"5d",x"5c",x"5b",x"5e"),
   579 => (x"4b",x"71",x"1e",x"0e"),
   580 => (x"73",x"4d",x"66",x"d4"),
   581 => (x"cc",x"c1",x"02",x"9b"),
   582 => (x"49",x"a3",x"c8",x"87"),
   583 => (x"c4",x"c1",x"02",x"69"),
   584 => (x"4c",x"a3",x"d0",x"87"),
   585 => (x"bf",x"ea",x"ec",x"c2"),
   586 => (x"6c",x"b9",x"ff",x"49"),
   587 => (x"d4",x"7e",x"99",x"4a"),
   588 => (x"cd",x"06",x"a9",x"66"),
   589 => (x"7c",x"7b",x"c0",x"87"),
   590 => (x"c4",x"4a",x"a3",x"cc"),
   591 => (x"79",x"6a",x"49",x"a3"),
   592 => (x"49",x"72",x"87",x"ca"),
   593 => (x"d4",x"99",x"c0",x"f8"),
   594 => (x"8d",x"71",x"4d",x"66"),
   595 => (x"29",x"c9",x"49",x"75"),
   596 => (x"49",x"73",x"1e",x"71"),
   597 => (x"c2",x"87",x"c7",x"fc"),
   598 => (x"73",x"1e",x"e6",x"e4"),
   599 => (x"87",x"d8",x"fd",x"49"),
   600 => (x"66",x"d4",x"86",x"c8"),
   601 => (x"e2",x"f6",x"26",x"7c"),
   602 => (x"5b",x"5e",x"0e",x"87"),
   603 => (x"f0",x"0e",x"5d",x"5c"),
   604 => (x"59",x"a6",x"d0",x"86"),
   605 => (x"4b",x"66",x"e4",x"c0"),
   606 => (x"ca",x"02",x"66",x"cc"),
   607 => (x"80",x"c8",x"48",x"87"),
   608 => (x"bf",x"6e",x"7e",x"70"),
   609 => (x"c0",x"87",x"c5",x"05"),
   610 => (x"87",x"ec",x"c3",x"48"),
   611 => (x"d0",x"4c",x"66",x"cc"),
   612 => (x"c4",x"49",x"73",x"84"),
   613 => (x"78",x"6c",x"48",x"a6"),
   614 => (x"c4",x"81",x"66",x"c4"),
   615 => (x"78",x"bf",x"6e",x"80"),
   616 => (x"06",x"a9",x"66",x"c8"),
   617 => (x"c4",x"49",x"87",x"c6"),
   618 => (x"4b",x"71",x"89",x"66"),
   619 => (x"01",x"ab",x"b7",x"c0"),
   620 => (x"c3",x"48",x"87",x"c4"),
   621 => (x"66",x"c4",x"87",x"c2"),
   622 => (x"98",x"ff",x"c7",x"48"),
   623 => (x"02",x"6e",x"7e",x"70"),
   624 => (x"c8",x"87",x"c9",x"c1"),
   625 => (x"89",x"6e",x"49",x"c0"),
   626 => (x"e4",x"c2",x"4a",x"71"),
   627 => (x"85",x"6e",x"4d",x"e6"),
   628 => (x"06",x"aa",x"b7",x"73"),
   629 => (x"72",x"4a",x"87",x"c1"),
   630 => (x"66",x"c4",x"48",x"49"),
   631 => (x"72",x"7c",x"70",x"80"),
   632 => (x"8a",x"c1",x"49",x"8b"),
   633 => (x"d9",x"02",x"99",x"71"),
   634 => (x"66",x"e0",x"c0",x"87"),
   635 => (x"c0",x"50",x"15",x"48"),
   636 => (x"c1",x"48",x"66",x"e0"),
   637 => (x"a6",x"e4",x"c0",x"80"),
   638 => (x"c1",x"49",x"72",x"58"),
   639 => (x"05",x"99",x"71",x"8a"),
   640 => (x"1e",x"c1",x"87",x"e7"),
   641 => (x"f9",x"49",x"66",x"d0"),
   642 => (x"86",x"c4",x"87",x"d4"),
   643 => (x"06",x"ab",x"b7",x"c0"),
   644 => (x"c0",x"87",x"e3",x"c1"),
   645 => (x"c7",x"4d",x"66",x"e0"),
   646 => (x"06",x"ab",x"b7",x"ff"),
   647 => (x"75",x"87",x"e2",x"c0"),
   648 => (x"49",x"66",x"d0",x"1e"),
   649 => (x"c8",x"87",x"d1",x"fa"),
   650 => (x"48",x"6c",x"85",x"c0"),
   651 => (x"70",x"80",x"c0",x"c8"),
   652 => (x"8b",x"c0",x"c8",x"7c"),
   653 => (x"66",x"d4",x"1e",x"c1"),
   654 => (x"87",x"e2",x"f8",x"49"),
   655 => (x"ee",x"c0",x"86",x"c8"),
   656 => (x"e6",x"e4",x"c2",x"87"),
   657 => (x"49",x"66",x"d0",x"1e"),
   658 => (x"c4",x"87",x"ed",x"f9"),
   659 => (x"e6",x"e4",x"c2",x"86"),
   660 => (x"48",x"49",x"73",x"4a"),
   661 => (x"7c",x"70",x"80",x"6c"),
   662 => (x"8b",x"c1",x"49",x"73"),
   663 => (x"ce",x"02",x"99",x"71"),
   664 => (x"7d",x"97",x"12",x"87"),
   665 => (x"49",x"73",x"85",x"c1"),
   666 => (x"99",x"71",x"8b",x"c1"),
   667 => (x"c0",x"87",x"f2",x"05"),
   668 => (x"fe",x"01",x"ab",x"b7"),
   669 => (x"48",x"c1",x"87",x"e1"),
   670 => (x"ce",x"f2",x"8e",x"f0"),
   671 => (x"5b",x"5e",x"0e",x"87"),
   672 => (x"71",x"0e",x"5d",x"5c"),
   673 => (x"c7",x"02",x"9b",x"4b"),
   674 => (x"4d",x"a3",x"c8",x"87"),
   675 => (x"87",x"c5",x"05",x"6d"),
   676 => (x"fd",x"c0",x"48",x"ff"),
   677 => (x"4c",x"a3",x"d0",x"87"),
   678 => (x"ff",x"c7",x"49",x"6c"),
   679 => (x"87",x"d8",x"05",x"99"),
   680 => (x"87",x"c9",x"02",x"6c"),
   681 => (x"49",x"73",x"1e",x"c1"),
   682 => (x"c4",x"87",x"f3",x"f6"),
   683 => (x"e6",x"e4",x"c2",x"86"),
   684 => (x"f8",x"49",x"73",x"1e"),
   685 => (x"86",x"c4",x"87",x"c2"),
   686 => (x"aa",x"6d",x"4a",x"6c"),
   687 => (x"ff",x"87",x"c4",x"04"),
   688 => (x"c1",x"87",x"cf",x"48"),
   689 => (x"49",x"72",x"7c",x"a2"),
   690 => (x"c2",x"99",x"ff",x"c7"),
   691 => (x"97",x"81",x"e6",x"e4"),
   692 => (x"f6",x"f0",x"48",x"69"),
   693 => (x"1e",x"73",x"1e",x"87"),
   694 => (x"02",x"9b",x"4b",x"71"),
   695 => (x"c2",x"87",x"e4",x"c0"),
   696 => (x"73",x"5b",x"d3",x"f1"),
   697 => (x"c2",x"8a",x"c2",x"4a"),
   698 => (x"49",x"bf",x"e6",x"ec"),
   699 => (x"ff",x"f0",x"c2",x"92"),
   700 => (x"80",x"72",x"48",x"bf"),
   701 => (x"58",x"d7",x"f1",x"c2"),
   702 => (x"30",x"c4",x"48",x"71"),
   703 => (x"58",x"f6",x"ec",x"c2"),
   704 => (x"c2",x"87",x"ed",x"c0"),
   705 => (x"c2",x"48",x"cf",x"f1"),
   706 => (x"78",x"bf",x"c3",x"f1"),
   707 => (x"48",x"d3",x"f1",x"c2"),
   708 => (x"bf",x"c7",x"f1",x"c2"),
   709 => (x"ee",x"ec",x"c2",x"78"),
   710 => (x"87",x"c9",x"02",x"bf"),
   711 => (x"bf",x"e6",x"ec",x"c2"),
   712 => (x"c7",x"31",x"c4",x"49"),
   713 => (x"cb",x"f1",x"c2",x"87"),
   714 => (x"31",x"c4",x"49",x"bf"),
   715 => (x"59",x"f6",x"ec",x"c2"),
   716 => (x"0e",x"87",x"dc",x"ef"),
   717 => (x"0e",x"5c",x"5b",x"5e"),
   718 => (x"4b",x"c0",x"4a",x"71"),
   719 => (x"c0",x"02",x"9a",x"72"),
   720 => (x"a2",x"da",x"87",x"e1"),
   721 => (x"4b",x"69",x"9f",x"49"),
   722 => (x"bf",x"ee",x"ec",x"c2"),
   723 => (x"d4",x"87",x"cf",x"02"),
   724 => (x"69",x"9f",x"49",x"a2"),
   725 => (x"ff",x"c0",x"4c",x"49"),
   726 => (x"34",x"d0",x"9c",x"ff"),
   727 => (x"4c",x"c0",x"87",x"c2"),
   728 => (x"73",x"b3",x"49",x"74"),
   729 => (x"87",x"ed",x"fd",x"49"),
   730 => (x"0e",x"87",x"e2",x"ee"),
   731 => (x"5d",x"5c",x"5b",x"5e"),
   732 => (x"71",x"86",x"f4",x"0e"),
   733 => (x"72",x"7e",x"c0",x"4a"),
   734 => (x"87",x"d8",x"02",x"9a"),
   735 => (x"48",x"e2",x"e4",x"c2"),
   736 => (x"e4",x"c2",x"78",x"c0"),
   737 => (x"f1",x"c2",x"48",x"da"),
   738 => (x"c2",x"78",x"bf",x"d3"),
   739 => (x"c2",x"48",x"de",x"e4"),
   740 => (x"78",x"bf",x"cf",x"f1"),
   741 => (x"48",x"c3",x"ed",x"c2"),
   742 => (x"ec",x"c2",x"50",x"c0"),
   743 => (x"c2",x"49",x"bf",x"f2"),
   744 => (x"4a",x"bf",x"e2",x"e4"),
   745 => (x"c4",x"03",x"aa",x"71"),
   746 => (x"49",x"72",x"87",x"ca"),
   747 => (x"c0",x"05",x"99",x"cf"),
   748 => (x"f5",x"c0",x"87",x"ea"),
   749 => (x"e4",x"c2",x"48",x"c7"),
   750 => (x"c2",x"78",x"bf",x"da"),
   751 => (x"c2",x"1e",x"e6",x"e4"),
   752 => (x"49",x"bf",x"da",x"e4"),
   753 => (x"48",x"da",x"e4",x"c2"),
   754 => (x"71",x"78",x"a1",x"c1"),
   755 => (x"87",x"fd",x"de",x"ff"),
   756 => (x"f5",x"c0",x"86",x"c4"),
   757 => (x"e4",x"c2",x"48",x"c3"),
   758 => (x"87",x"cc",x"78",x"e6"),
   759 => (x"bf",x"c3",x"f5",x"c0"),
   760 => (x"80",x"e0",x"c0",x"48"),
   761 => (x"58",x"c7",x"f5",x"c0"),
   762 => (x"bf",x"e2",x"e4",x"c2"),
   763 => (x"c2",x"80",x"c1",x"48"),
   764 => (x"27",x"58",x"e6",x"e4"),
   765 => (x"00",x"00",x"0d",x"43"),
   766 => (x"4d",x"bf",x"97",x"bf"),
   767 => (x"e3",x"c2",x"02",x"9d"),
   768 => (x"ad",x"e5",x"c3",x"87"),
   769 => (x"87",x"dc",x"c2",x"02"),
   770 => (x"bf",x"c3",x"f5",x"c0"),
   771 => (x"49",x"a3",x"cb",x"4b"),
   772 => (x"ac",x"cf",x"4c",x"11"),
   773 => (x"87",x"d2",x"c1",x"05"),
   774 => (x"99",x"df",x"49",x"75"),
   775 => (x"91",x"cd",x"89",x"c1"),
   776 => (x"81",x"f6",x"ec",x"c2"),
   777 => (x"12",x"4a",x"a3",x"c1"),
   778 => (x"4a",x"a3",x"c3",x"51"),
   779 => (x"a3",x"c5",x"51",x"12"),
   780 => (x"c7",x"51",x"12",x"4a"),
   781 => (x"51",x"12",x"4a",x"a3"),
   782 => (x"12",x"4a",x"a3",x"c9"),
   783 => (x"4a",x"a3",x"ce",x"51"),
   784 => (x"a3",x"d0",x"51",x"12"),
   785 => (x"d2",x"51",x"12",x"4a"),
   786 => (x"51",x"12",x"4a",x"a3"),
   787 => (x"12",x"4a",x"a3",x"d4"),
   788 => (x"4a",x"a3",x"d6",x"51"),
   789 => (x"a3",x"d8",x"51",x"12"),
   790 => (x"dc",x"51",x"12",x"4a"),
   791 => (x"51",x"12",x"4a",x"a3"),
   792 => (x"12",x"4a",x"a3",x"de"),
   793 => (x"c0",x"7e",x"c1",x"51"),
   794 => (x"49",x"74",x"87",x"fa"),
   795 => (x"c0",x"05",x"99",x"c8"),
   796 => (x"49",x"74",x"87",x"eb"),
   797 => (x"d1",x"05",x"99",x"d0"),
   798 => (x"02",x"66",x"dc",x"87"),
   799 => (x"73",x"87",x"cb",x"c0"),
   800 => (x"0f",x"66",x"dc",x"49"),
   801 => (x"c0",x"02",x"98",x"70"),
   802 => (x"05",x"6e",x"87",x"d3"),
   803 => (x"c2",x"87",x"c6",x"c0"),
   804 => (x"c0",x"48",x"f6",x"ec"),
   805 => (x"c3",x"f5",x"c0",x"50"),
   806 => (x"e1",x"c2",x"48",x"bf"),
   807 => (x"c3",x"ed",x"c2",x"87"),
   808 => (x"7e",x"50",x"c0",x"48"),
   809 => (x"bf",x"f2",x"ec",x"c2"),
   810 => (x"e2",x"e4",x"c2",x"49"),
   811 => (x"aa",x"71",x"4a",x"bf"),
   812 => (x"87",x"f6",x"fb",x"04"),
   813 => (x"bf",x"d3",x"f1",x"c2"),
   814 => (x"87",x"c8",x"c0",x"05"),
   815 => (x"bf",x"ee",x"ec",x"c2"),
   816 => (x"87",x"f8",x"c1",x"02"),
   817 => (x"bf",x"de",x"e4",x"c2"),
   818 => (x"87",x"c7",x"e9",x"49"),
   819 => (x"e4",x"c2",x"49",x"70"),
   820 => (x"a6",x"c4",x"59",x"e2"),
   821 => (x"de",x"e4",x"c2",x"48"),
   822 => (x"ec",x"c2",x"78",x"bf"),
   823 => (x"c0",x"02",x"bf",x"ee"),
   824 => (x"66",x"c4",x"87",x"d8"),
   825 => (x"ff",x"ff",x"cf",x"49"),
   826 => (x"a9",x"99",x"f8",x"ff"),
   827 => (x"87",x"c5",x"c0",x"02"),
   828 => (x"e1",x"c0",x"4c",x"c0"),
   829 => (x"c0",x"4c",x"c1",x"87"),
   830 => (x"66",x"c4",x"87",x"dc"),
   831 => (x"f8",x"ff",x"cf",x"49"),
   832 => (x"c0",x"02",x"a9",x"99"),
   833 => (x"a6",x"c8",x"87",x"c8"),
   834 => (x"c0",x"78",x"c0",x"48"),
   835 => (x"a6",x"c8",x"87",x"c5"),
   836 => (x"c8",x"78",x"c1",x"48"),
   837 => (x"9c",x"74",x"4c",x"66"),
   838 => (x"87",x"e0",x"c0",x"05"),
   839 => (x"c2",x"49",x"66",x"c4"),
   840 => (x"e6",x"ec",x"c2",x"89"),
   841 => (x"c2",x"91",x"4a",x"bf"),
   842 => (x"4a",x"bf",x"ff",x"f0"),
   843 => (x"48",x"da",x"e4",x"c2"),
   844 => (x"c2",x"78",x"a1",x"72"),
   845 => (x"c0",x"48",x"e2",x"e4"),
   846 => (x"87",x"de",x"f9",x"78"),
   847 => (x"8e",x"f4",x"48",x"c0"),
   848 => (x"00",x"87",x"c8",x"e7"),
   849 => (x"ff",x"00",x"00",x"00"),
   850 => (x"53",x"ff",x"ff",x"ff"),
   851 => (x"5c",x"00",x"00",x"0d"),
   852 => (x"46",x"00",x"00",x"0d"),
   853 => (x"32",x"33",x"54",x"41"),
   854 => (x"00",x"20",x"20",x"20"),
   855 => (x"31",x"54",x"41",x"46"),
   856 => (x"20",x"20",x"20",x"36"),
   857 => (x"f1",x"c2",x"1e",x"00"),
   858 => (x"dd",x"48",x"bf",x"d8"),
   859 => (x"87",x"c9",x"05",x"a8"),
   860 => (x"87",x"cd",x"c2",x"c1"),
   861 => (x"c8",x"4a",x"49",x"70"),
   862 => (x"48",x"d4",x"ff",x"87"),
   863 => (x"68",x"78",x"ff",x"c3"),
   864 => (x"26",x"48",x"72",x"4a"),
   865 => (x"f1",x"c2",x"1e",x"4f"),
   866 => (x"dd",x"48",x"bf",x"d8"),
   867 => (x"87",x"c6",x"05",x"a8"),
   868 => (x"87",x"d9",x"c1",x"c1"),
   869 => (x"d4",x"ff",x"87",x"d9"),
   870 => (x"78",x"ff",x"c3",x"48"),
   871 => (x"c0",x"48",x"d0",x"ff"),
   872 => (x"d4",x"ff",x"78",x"e1"),
   873 => (x"c2",x"78",x"d4",x"48"),
   874 => (x"ff",x"48",x"d7",x"f1"),
   875 => (x"26",x"50",x"bf",x"d4"),
   876 => (x"d0",x"ff",x"1e",x"4f"),
   877 => (x"78",x"e0",x"c0",x"48"),
   878 => (x"fe",x"1e",x"4f",x"26"),
   879 => (x"49",x"70",x"87",x"e7"),
   880 => (x"87",x"c6",x"02",x"99"),
   881 => (x"05",x"a9",x"fb",x"c0"),
   882 => (x"48",x"71",x"87",x"f1"),
   883 => (x"5e",x"0e",x"4f",x"26"),
   884 => (x"71",x"0e",x"5c",x"5b"),
   885 => (x"fe",x"4c",x"c0",x"4b"),
   886 => (x"49",x"70",x"87",x"cb"),
   887 => (x"f9",x"c0",x"02",x"99"),
   888 => (x"a9",x"ec",x"c0",x"87"),
   889 => (x"87",x"f2",x"c0",x"02"),
   890 => (x"02",x"a9",x"fb",x"c0"),
   891 => (x"cc",x"87",x"eb",x"c0"),
   892 => (x"03",x"ac",x"b7",x"66"),
   893 => (x"66",x"d0",x"87",x"c7"),
   894 => (x"71",x"87",x"c2",x"02"),
   895 => (x"02",x"99",x"71",x"53"),
   896 => (x"84",x"c1",x"87",x"c2"),
   897 => (x"70",x"87",x"de",x"fd"),
   898 => (x"cd",x"02",x"99",x"49"),
   899 => (x"a9",x"ec",x"c0",x"87"),
   900 => (x"c0",x"87",x"c7",x"02"),
   901 => (x"ff",x"05",x"a9",x"fb"),
   902 => (x"66",x"d0",x"87",x"d5"),
   903 => (x"c0",x"87",x"c3",x"02"),
   904 => (x"ec",x"c0",x"7b",x"97"),
   905 => (x"87",x"c4",x"05",x"a9"),
   906 => (x"87",x"c5",x"4a",x"74"),
   907 => (x"0a",x"c0",x"4a",x"74"),
   908 => (x"c2",x"48",x"72",x"8a"),
   909 => (x"26",x"4d",x"26",x"87"),
   910 => (x"26",x"4b",x"26",x"4c"),
   911 => (x"e4",x"fc",x"1e",x"4f"),
   912 => (x"4a",x"49",x"70",x"87"),
   913 => (x"04",x"aa",x"f0",x"c0"),
   914 => (x"f9",x"c0",x"87",x"c9"),
   915 => (x"87",x"c3",x"01",x"aa"),
   916 => (x"c1",x"8a",x"f0",x"c0"),
   917 => (x"c9",x"04",x"aa",x"c1"),
   918 => (x"aa",x"da",x"c1",x"87"),
   919 => (x"c0",x"87",x"c3",x"01"),
   920 => (x"48",x"72",x"8a",x"f7"),
   921 => (x"5e",x"0e",x"4f",x"26"),
   922 => (x"71",x"0e",x"5c",x"5b"),
   923 => (x"4c",x"d4",x"ff",x"4a"),
   924 => (x"e9",x"c0",x"49",x"72"),
   925 => (x"9b",x"4b",x"70",x"87"),
   926 => (x"c1",x"87",x"c2",x"02"),
   927 => (x"48",x"d0",x"ff",x"8b"),
   928 => (x"d5",x"c1",x"78",x"c5"),
   929 => (x"c6",x"49",x"73",x"7c"),
   930 => (x"c3",x"e7",x"c1",x"31"),
   931 => (x"48",x"4a",x"bf",x"97"),
   932 => (x"7c",x"70",x"b0",x"71"),
   933 => (x"c4",x"48",x"d0",x"ff"),
   934 => (x"fe",x"48",x"73",x"78"),
   935 => (x"5e",x"0e",x"87",x"d9"),
   936 => (x"0e",x"5d",x"5c",x"5b"),
   937 => (x"4b",x"71",x"86",x"f8"),
   938 => (x"fe",x"c0",x"7e",x"c0"),
   939 => (x"49",x"bf",x"97",x"c4"),
   940 => (x"ee",x"c0",x"05",x"99"),
   941 => (x"49",x"a3",x"c8",x"87"),
   942 => (x"c1",x"49",x"69",x"97"),
   943 => (x"dd",x"05",x"a9",x"c1"),
   944 => (x"49",x"a3",x"c9",x"87"),
   945 => (x"c1",x"49",x"69",x"97"),
   946 => (x"d1",x"05",x"a9",x"d2"),
   947 => (x"49",x"a3",x"ca",x"87"),
   948 => (x"c1",x"49",x"69",x"97"),
   949 => (x"c5",x"05",x"a9",x"c3"),
   950 => (x"c2",x"48",x"df",x"87"),
   951 => (x"48",x"c0",x"87",x"e1"),
   952 => (x"fa",x"87",x"dc",x"c2"),
   953 => (x"4c",x"c0",x"87",x"df"),
   954 => (x"97",x"c4",x"fe",x"c0"),
   955 => (x"a9",x"c0",x"49",x"bf"),
   956 => (x"fb",x"87",x"cf",x"04"),
   957 => (x"84",x"c1",x"87",x"c4"),
   958 => (x"97",x"c4",x"fe",x"c0"),
   959 => (x"06",x"ac",x"49",x"bf"),
   960 => (x"fe",x"c0",x"87",x"f1"),
   961 => (x"02",x"bf",x"97",x"c4"),
   962 => (x"d8",x"f9",x"87",x"cf"),
   963 => (x"99",x"49",x"70",x"87"),
   964 => (x"c0",x"87",x"c6",x"02"),
   965 => (x"f1",x"05",x"a9",x"ec"),
   966 => (x"f9",x"4c",x"c0",x"87"),
   967 => (x"4d",x"70",x"87",x"c7"),
   968 => (x"c8",x"87",x"c2",x"f9"),
   969 => (x"fc",x"f8",x"58",x"a6"),
   970 => (x"c1",x"4a",x"70",x"87"),
   971 => (x"49",x"a3",x"c8",x"84"),
   972 => (x"ad",x"49",x"69",x"97"),
   973 => (x"c0",x"87",x"c7",x"02"),
   974 => (x"c0",x"05",x"ad",x"ff"),
   975 => (x"a3",x"c9",x"87",x"e7"),
   976 => (x"49",x"69",x"97",x"49"),
   977 => (x"02",x"a9",x"66",x"c4"),
   978 => (x"c0",x"48",x"87",x"c7"),
   979 => (x"d4",x"05",x"a8",x"ff"),
   980 => (x"49",x"a3",x"ca",x"87"),
   981 => (x"aa",x"49",x"69",x"97"),
   982 => (x"c0",x"87",x"c6",x"02"),
   983 => (x"c4",x"05",x"aa",x"ff"),
   984 => (x"d0",x"7e",x"c1",x"87"),
   985 => (x"ad",x"ec",x"c0",x"87"),
   986 => (x"c0",x"87",x"c6",x"02"),
   987 => (x"c4",x"05",x"ad",x"fb"),
   988 => (x"c1",x"4c",x"c0",x"87"),
   989 => (x"fe",x"02",x"6e",x"7e"),
   990 => (x"f4",x"f8",x"87",x"e1"),
   991 => (x"f8",x"48",x"74",x"87"),
   992 => (x"87",x"f1",x"fa",x"8e"),
   993 => (x"5b",x"5e",x"0e",x"00"),
   994 => (x"f8",x"0e",x"5d",x"5c"),
   995 => (x"ff",x"4d",x"71",x"86"),
   996 => (x"1e",x"75",x"4b",x"d4"),
   997 => (x"49",x"dc",x"f1",x"c2"),
   998 => (x"87",x"e9",x"df",x"ff"),
   999 => (x"98",x"70",x"86",x"c4"),
  1000 => (x"87",x"fb",x"c4",x"02"),
  1001 => (x"bf",x"c5",x"e7",x"c1"),
  1002 => (x"fa",x"49",x"75",x"7e"),
  1003 => (x"a8",x"de",x"87",x"f8"),
  1004 => (x"87",x"eb",x"c0",x"05"),
  1005 => (x"f6",x"c0",x"49",x"75"),
  1006 => (x"98",x"70",x"87",x"e5"),
  1007 => (x"c2",x"87",x"db",x"02"),
  1008 => (x"1e",x"bf",x"c0",x"f6"),
  1009 => (x"c0",x"49",x"e1",x"c0"),
  1010 => (x"c4",x"87",x"f4",x"f3"),
  1011 => (x"c3",x"e7",x"c1",x"86"),
  1012 => (x"c2",x"50",x"c0",x"48"),
  1013 => (x"fe",x"49",x"cc",x"f6"),
  1014 => (x"48",x"c1",x"87",x"eb"),
  1015 => (x"ff",x"87",x"c2",x"c4"),
  1016 => (x"78",x"c5",x"48",x"d0"),
  1017 => (x"c0",x"7b",x"d6",x"c1"),
  1018 => (x"49",x"a2",x"75",x"4a"),
  1019 => (x"82",x"c1",x"7b",x"11"),
  1020 => (x"04",x"aa",x"b7",x"cb"),
  1021 => (x"4a",x"cc",x"87",x"f3"),
  1022 => (x"c1",x"7b",x"ff",x"c3"),
  1023 => (x"b7",x"e0",x"c0",x"82"),
  1024 => (x"87",x"f4",x"04",x"aa"),
  1025 => (x"c4",x"48",x"d0",x"ff"),
  1026 => (x"7b",x"ff",x"c3",x"78"),
  1027 => (x"d3",x"c1",x"78",x"c5"),
  1028 => (x"c4",x"7b",x"c1",x"7b"),
  1029 => (x"c0",x"48",x"6e",x"78"),
  1030 => (x"c2",x"06",x"a8",x"b7"),
  1031 => (x"f1",x"c2",x"87",x"f0"),
  1032 => (x"6e",x"4c",x"bf",x"e4"),
  1033 => (x"70",x"88",x"74",x"48"),
  1034 => (x"02",x"9c",x"74",x"7e"),
  1035 => (x"c2",x"87",x"fd",x"c1"),
  1036 => (x"c4",x"4d",x"e6",x"e4"),
  1037 => (x"c0",x"c8",x"48",x"a6"),
  1038 => (x"b7",x"c0",x"8c",x"78"),
  1039 => (x"87",x"c6",x"03",x"ac"),
  1040 => (x"78",x"a4",x"c0",x"c8"),
  1041 => (x"f1",x"c2",x"4c",x"c0"),
  1042 => (x"49",x"bf",x"97",x"d7"),
  1043 => (x"d1",x"02",x"99",x"d0"),
  1044 => (x"c2",x"1e",x"c0",x"87"),
  1045 => (x"e1",x"49",x"dc",x"f1"),
  1046 => (x"86",x"c4",x"87",x"de"),
  1047 => (x"c0",x"4a",x"49",x"70"),
  1048 => (x"e4",x"c2",x"87",x"ee"),
  1049 => (x"f1",x"c2",x"1e",x"e6"),
  1050 => (x"cb",x"e1",x"49",x"dc"),
  1051 => (x"70",x"86",x"c4",x"87"),
  1052 => (x"d0",x"ff",x"4a",x"49"),
  1053 => (x"78",x"c5",x"c8",x"48"),
  1054 => (x"15",x"7b",x"d4",x"c1"),
  1055 => (x"48",x"66",x"c4",x"7b"),
  1056 => (x"a6",x"c8",x"88",x"c1"),
  1057 => (x"05",x"98",x"70",x"58"),
  1058 => (x"ff",x"87",x"f0",x"ff"),
  1059 => (x"78",x"c4",x"48",x"d0"),
  1060 => (x"c5",x"05",x"9a",x"72"),
  1061 => (x"c1",x"48",x"c0",x"87"),
  1062 => (x"1e",x"c1",x"87",x"c7"),
  1063 => (x"49",x"dc",x"f1",x"c2"),
  1064 => (x"87",x"fa",x"de",x"ff"),
  1065 => (x"9c",x"74",x"86",x"c4"),
  1066 => (x"87",x"c3",x"fe",x"05"),
  1067 => (x"b7",x"c0",x"48",x"6e"),
  1068 => (x"87",x"d1",x"06",x"a8"),
  1069 => (x"48",x"dc",x"f1",x"c2"),
  1070 => (x"80",x"d0",x"78",x"c0"),
  1071 => (x"80",x"f4",x"78",x"c0"),
  1072 => (x"bf",x"e8",x"f1",x"c2"),
  1073 => (x"c0",x"48",x"6e",x"78"),
  1074 => (x"fd",x"01",x"a8",x"b7"),
  1075 => (x"d0",x"ff",x"87",x"d0"),
  1076 => (x"c1",x"78",x"c5",x"48"),
  1077 => (x"7b",x"c0",x"7b",x"d3"),
  1078 => (x"48",x"c1",x"78",x"c4"),
  1079 => (x"c0",x"87",x"c2",x"c0"),
  1080 => (x"26",x"8e",x"f8",x"48"),
  1081 => (x"26",x"4c",x"26",x"4d"),
  1082 => (x"0e",x"4f",x"26",x"4b"),
  1083 => (x"5d",x"5c",x"5b",x"5e"),
  1084 => (x"4b",x"71",x"1e",x"0e"),
  1085 => (x"ab",x"4d",x"4c",x"c0"),
  1086 => (x"87",x"e8",x"c0",x"04"),
  1087 => (x"1e",x"de",x"fa",x"c0"),
  1088 => (x"c4",x"02",x"9d",x"75"),
  1089 => (x"c2",x"4a",x"c0",x"87"),
  1090 => (x"72",x"4a",x"c1",x"87"),
  1091 => (x"87",x"db",x"e9",x"49"),
  1092 => (x"7e",x"70",x"86",x"c4"),
  1093 => (x"05",x"6e",x"84",x"c1"),
  1094 => (x"4c",x"73",x"87",x"c2"),
  1095 => (x"ac",x"73",x"85",x"c1"),
  1096 => (x"87",x"d8",x"ff",x"06"),
  1097 => (x"fe",x"26",x"48",x"6e"),
  1098 => (x"71",x"1e",x"87",x"f9"),
  1099 => (x"05",x"66",x"c4",x"4a"),
  1100 => (x"49",x"72",x"87",x"c5"),
  1101 => (x"26",x"87",x"ce",x"f9"),
  1102 => (x"5b",x"5e",x"0e",x"4f"),
  1103 => (x"1e",x"0e",x"5d",x"5c"),
  1104 => (x"de",x"49",x"4c",x"71"),
  1105 => (x"c4",x"f2",x"c2",x"91"),
  1106 => (x"97",x"85",x"71",x"4d"),
  1107 => (x"dc",x"c1",x"02",x"6d"),
  1108 => (x"f0",x"f1",x"c2",x"87"),
  1109 => (x"82",x"74",x"4a",x"bf"),
  1110 => (x"ce",x"fe",x"49",x"72"),
  1111 => (x"6e",x"7e",x"70",x"87"),
  1112 => (x"87",x"f2",x"c0",x"02"),
  1113 => (x"4b",x"f8",x"f1",x"c2"),
  1114 => (x"49",x"cb",x"4a",x"6e"),
  1115 => (x"87",x"f8",x"fc",x"fe"),
  1116 => (x"93",x"cb",x"4b",x"74"),
  1117 => (x"83",x"d7",x"e7",x"c1"),
  1118 => (x"c6",x"c1",x"83",x"c4"),
  1119 => (x"49",x"74",x"7b",x"f1"),
  1120 => (x"87",x"fc",x"ca",x"c1"),
  1121 => (x"e7",x"c1",x"7b",x"75"),
  1122 => (x"49",x"bf",x"97",x"c4"),
  1123 => (x"f8",x"f1",x"c2",x"1e"),
  1124 => (x"87",x"d6",x"fe",x"49"),
  1125 => (x"49",x"74",x"86",x"c4"),
  1126 => (x"87",x"e4",x"ca",x"c1"),
  1127 => (x"cc",x"c1",x"49",x"c0"),
  1128 => (x"f1",x"c2",x"87",x"c3"),
  1129 => (x"78",x"c0",x"48",x"d8"),
  1130 => (x"d9",x"dd",x"49",x"c1"),
  1131 => (x"f2",x"fc",x"26",x"87"),
  1132 => (x"61",x"6f",x"4c",x"87"),
  1133 => (x"67",x"6e",x"69",x"64"),
  1134 => (x"00",x"2e",x"2e",x"2e"),
  1135 => (x"5c",x"5b",x"5e",x"0e"),
  1136 => (x"4a",x"4b",x"71",x"0e"),
  1137 => (x"bf",x"f0",x"f1",x"c2"),
  1138 => (x"fc",x"49",x"72",x"82"),
  1139 => (x"4c",x"70",x"87",x"dd"),
  1140 => (x"87",x"c4",x"02",x"9c"),
  1141 => (x"87",x"db",x"e5",x"49"),
  1142 => (x"48",x"f0",x"f1",x"c2"),
  1143 => (x"49",x"c1",x"78",x"c0"),
  1144 => (x"fb",x"87",x"e3",x"dc"),
  1145 => (x"5e",x"0e",x"87",x"ff"),
  1146 => (x"0e",x"5d",x"5c",x"5b"),
  1147 => (x"e4",x"c2",x"86",x"f4"),
  1148 => (x"4c",x"c0",x"4d",x"e6"),
  1149 => (x"c0",x"48",x"a6",x"c4"),
  1150 => (x"f0",x"f1",x"c2",x"78"),
  1151 => (x"a9",x"c0",x"49",x"bf"),
  1152 => (x"87",x"c1",x"c1",x"06"),
  1153 => (x"48",x"e6",x"e4",x"c2"),
  1154 => (x"f8",x"c0",x"02",x"98"),
  1155 => (x"de",x"fa",x"c0",x"87"),
  1156 => (x"02",x"66",x"c8",x"1e"),
  1157 => (x"a6",x"c4",x"87",x"c7"),
  1158 => (x"c5",x"78",x"c0",x"48"),
  1159 => (x"48",x"a6",x"c4",x"87"),
  1160 => (x"66",x"c4",x"78",x"c1"),
  1161 => (x"87",x"c3",x"e5",x"49"),
  1162 => (x"4d",x"70",x"86",x"c4"),
  1163 => (x"66",x"c4",x"84",x"c1"),
  1164 => (x"c8",x"80",x"c1",x"48"),
  1165 => (x"f1",x"c2",x"58",x"a6"),
  1166 => (x"ac",x"49",x"bf",x"f0"),
  1167 => (x"75",x"87",x"c6",x"03"),
  1168 => (x"c8",x"ff",x"05",x"9d"),
  1169 => (x"75",x"4c",x"c0",x"87"),
  1170 => (x"e0",x"c3",x"02",x"9d"),
  1171 => (x"de",x"fa",x"c0",x"87"),
  1172 => (x"02",x"66",x"c8",x"1e"),
  1173 => (x"a6",x"cc",x"87",x"c7"),
  1174 => (x"c5",x"78",x"c0",x"48"),
  1175 => (x"48",x"a6",x"cc",x"87"),
  1176 => (x"66",x"cc",x"78",x"c1"),
  1177 => (x"87",x"c3",x"e4",x"49"),
  1178 => (x"7e",x"70",x"86",x"c4"),
  1179 => (x"e9",x"c2",x"02",x"6e"),
  1180 => (x"cb",x"49",x"6e",x"87"),
  1181 => (x"49",x"69",x"97",x"81"),
  1182 => (x"c1",x"02",x"99",x"d0"),
  1183 => (x"c6",x"c1",x"87",x"d6"),
  1184 => (x"49",x"74",x"4a",x"fc"),
  1185 => (x"e7",x"c1",x"91",x"cb"),
  1186 => (x"79",x"72",x"81",x"d7"),
  1187 => (x"ff",x"c3",x"81",x"c8"),
  1188 => (x"de",x"49",x"74",x"51"),
  1189 => (x"c4",x"f2",x"c2",x"91"),
  1190 => (x"c2",x"85",x"71",x"4d"),
  1191 => (x"c1",x"7d",x"97",x"c1"),
  1192 => (x"e0",x"c0",x"49",x"a5"),
  1193 => (x"f6",x"ec",x"c2",x"51"),
  1194 => (x"d2",x"02",x"bf",x"97"),
  1195 => (x"c2",x"84",x"c1",x"87"),
  1196 => (x"ec",x"c2",x"4b",x"a5"),
  1197 => (x"49",x"db",x"4a",x"f6"),
  1198 => (x"87",x"ec",x"f7",x"fe"),
  1199 => (x"cd",x"87",x"db",x"c1"),
  1200 => (x"51",x"c0",x"49",x"a5"),
  1201 => (x"a5",x"c2",x"84",x"c1"),
  1202 => (x"cb",x"4a",x"6e",x"4b"),
  1203 => (x"d7",x"f7",x"fe",x"49"),
  1204 => (x"87",x"c6",x"c1",x"87"),
  1205 => (x"4a",x"f9",x"c4",x"c1"),
  1206 => (x"91",x"cb",x"49",x"74"),
  1207 => (x"81",x"d7",x"e7",x"c1"),
  1208 => (x"ec",x"c2",x"79",x"72"),
  1209 => (x"02",x"bf",x"97",x"f6"),
  1210 => (x"49",x"74",x"87",x"d8"),
  1211 => (x"84",x"c1",x"91",x"de"),
  1212 => (x"4b",x"c4",x"f2",x"c2"),
  1213 => (x"ec",x"c2",x"83",x"71"),
  1214 => (x"49",x"dd",x"4a",x"f6"),
  1215 => (x"87",x"e8",x"f6",x"fe"),
  1216 => (x"4b",x"74",x"87",x"d8"),
  1217 => (x"f2",x"c2",x"93",x"de"),
  1218 => (x"a3",x"cb",x"83",x"c4"),
  1219 => (x"c1",x"51",x"c0",x"49"),
  1220 => (x"4a",x"6e",x"73",x"84"),
  1221 => (x"f6",x"fe",x"49",x"cb"),
  1222 => (x"66",x"c4",x"87",x"ce"),
  1223 => (x"c8",x"80",x"c1",x"48"),
  1224 => (x"ac",x"c7",x"58",x"a6"),
  1225 => (x"87",x"c5",x"c0",x"03"),
  1226 => (x"e0",x"fc",x"05",x"6e"),
  1227 => (x"f4",x"48",x"74",x"87"),
  1228 => (x"87",x"ef",x"f6",x"8e"),
  1229 => (x"71",x"1e",x"73",x"1e"),
  1230 => (x"91",x"cb",x"49",x"4b"),
  1231 => (x"81",x"d7",x"e7",x"c1"),
  1232 => (x"c1",x"4a",x"a1",x"c8"),
  1233 => (x"12",x"48",x"c3",x"e7"),
  1234 => (x"4a",x"a1",x"c9",x"50"),
  1235 => (x"48",x"c4",x"fe",x"c0"),
  1236 => (x"81",x"ca",x"50",x"12"),
  1237 => (x"48",x"c4",x"e7",x"c1"),
  1238 => (x"e7",x"c1",x"50",x"11"),
  1239 => (x"49",x"bf",x"97",x"c4"),
  1240 => (x"f7",x"49",x"c0",x"1e"),
  1241 => (x"f1",x"c2",x"87",x"c4"),
  1242 => (x"78",x"de",x"48",x"d8"),
  1243 => (x"d5",x"d6",x"49",x"c1"),
  1244 => (x"f2",x"f5",x"26",x"87"),
  1245 => (x"4a",x"71",x"1e",x"87"),
  1246 => (x"c1",x"91",x"cb",x"49"),
  1247 => (x"c8",x"81",x"d7",x"e7"),
  1248 => (x"c2",x"48",x"11",x"81"),
  1249 => (x"c2",x"58",x"dc",x"f1"),
  1250 => (x"c0",x"48",x"f0",x"f1"),
  1251 => (x"d5",x"49",x"c1",x"78"),
  1252 => (x"4f",x"26",x"87",x"f4"),
  1253 => (x"c1",x"49",x"c0",x"1e"),
  1254 => (x"26",x"87",x"ca",x"c4"),
  1255 => (x"99",x"71",x"1e",x"4f"),
  1256 => (x"c1",x"87",x"d2",x"02"),
  1257 => (x"c0",x"48",x"ec",x"e8"),
  1258 => (x"c1",x"80",x"f7",x"50"),
  1259 => (x"c1",x"40",x"f5",x"cd"),
  1260 => (x"ce",x"78",x"d0",x"e7"),
  1261 => (x"e8",x"e8",x"c1",x"87"),
  1262 => (x"c9",x"e7",x"c1",x"48"),
  1263 => (x"c1",x"80",x"fc",x"78"),
  1264 => (x"26",x"78",x"d4",x"ce"),
  1265 => (x"5b",x"5e",x"0e",x"4f"),
  1266 => (x"4c",x"71",x"0e",x"5c"),
  1267 => (x"c1",x"92",x"cb",x"4a"),
  1268 => (x"c8",x"82",x"d7",x"e7"),
  1269 => (x"a2",x"c9",x"49",x"a2"),
  1270 => (x"4b",x"6b",x"97",x"4b"),
  1271 => (x"49",x"69",x"97",x"1e"),
  1272 => (x"12",x"82",x"ca",x"1e"),
  1273 => (x"f6",x"e4",x"c0",x"49"),
  1274 => (x"d4",x"49",x"c0",x"87"),
  1275 => (x"49",x"74",x"87",x"d8"),
  1276 => (x"87",x"cc",x"c1",x"c1"),
  1277 => (x"ec",x"f3",x"8e",x"f8"),
  1278 => (x"1e",x"73",x"1e",x"87"),
  1279 => (x"ff",x"49",x"4b",x"71"),
  1280 => (x"49",x"73",x"87",x"c3"),
  1281 => (x"f3",x"87",x"fe",x"fe"),
  1282 => (x"73",x"1e",x"87",x"dd"),
  1283 => (x"c6",x"4b",x"71",x"1e"),
  1284 => (x"db",x"02",x"4a",x"a3"),
  1285 => (x"02",x"8a",x"c1",x"87"),
  1286 => (x"02",x"8a",x"87",x"d6"),
  1287 => (x"8a",x"87",x"da",x"c1"),
  1288 => (x"87",x"fc",x"c0",x"02"),
  1289 => (x"e1",x"c0",x"02",x"8a"),
  1290 => (x"cb",x"02",x"8a",x"87"),
  1291 => (x"87",x"db",x"c1",x"87"),
  1292 => (x"c0",x"fd",x"49",x"c7"),
  1293 => (x"87",x"de",x"c1",x"87"),
  1294 => (x"bf",x"f0",x"f1",x"c2"),
  1295 => (x"87",x"cb",x"c1",x"02"),
  1296 => (x"c2",x"88",x"c1",x"48"),
  1297 => (x"c1",x"58",x"f4",x"f1"),
  1298 => (x"f1",x"c2",x"87",x"c1"),
  1299 => (x"c0",x"02",x"bf",x"f4"),
  1300 => (x"f1",x"c2",x"87",x"f9"),
  1301 => (x"c1",x"48",x"bf",x"f0"),
  1302 => (x"f4",x"f1",x"c2",x"80"),
  1303 => (x"87",x"eb",x"c0",x"58"),
  1304 => (x"bf",x"f0",x"f1",x"c2"),
  1305 => (x"c2",x"89",x"c6",x"49"),
  1306 => (x"c0",x"59",x"f4",x"f1"),
  1307 => (x"da",x"03",x"a9",x"b7"),
  1308 => (x"f0",x"f1",x"c2",x"87"),
  1309 => (x"d2",x"78",x"c0",x"48"),
  1310 => (x"f4",x"f1",x"c2",x"87"),
  1311 => (x"87",x"cb",x"02",x"bf"),
  1312 => (x"bf",x"f0",x"f1",x"c2"),
  1313 => (x"c2",x"80",x"c6",x"48"),
  1314 => (x"c0",x"58",x"f4",x"f1"),
  1315 => (x"87",x"f6",x"d1",x"49"),
  1316 => (x"fe",x"c0",x"49",x"73"),
  1317 => (x"ce",x"f1",x"87",x"ea"),
  1318 => (x"1e",x"73",x"1e",x"87"),
  1319 => (x"f1",x"c2",x"4b",x"71"),
  1320 => (x"78",x"dd",x"48",x"d8"),
  1321 => (x"dd",x"d1",x"49",x"c0"),
  1322 => (x"c0",x"49",x"73",x"87"),
  1323 => (x"f0",x"87",x"d1",x"fe"),
  1324 => (x"5e",x"0e",x"87",x"f5"),
  1325 => (x"0e",x"5d",x"5c",x"5b"),
  1326 => (x"d8",x"86",x"cc",x"ff"),
  1327 => (x"a6",x"c8",x"59",x"a6"),
  1328 => (x"c4",x"78",x"c0",x"48"),
  1329 => (x"66",x"c8",x"c1",x"80"),
  1330 => (x"c1",x"80",x"c4",x"78"),
  1331 => (x"f4",x"f1",x"c2",x"78"),
  1332 => (x"c2",x"78",x"c1",x"48"),
  1333 => (x"48",x"bf",x"d8",x"f1"),
  1334 => (x"cb",x"05",x"a8",x"de"),
  1335 => (x"87",x"c6",x"f4",x"87"),
  1336 => (x"a6",x"cc",x"49",x"70"),
  1337 => (x"87",x"d0",x"cf",x"59"),
  1338 => (x"e3",x"87",x"da",x"e2"),
  1339 => (x"f4",x"e1",x"87",x"cc"),
  1340 => (x"d4",x"4c",x"70",x"87"),
  1341 => (x"fc",x"c1",x"05",x"66"),
  1342 => (x"66",x"c4",x"c1",x"87"),
  1343 => (x"70",x"80",x"c4",x"48"),
  1344 => (x"48",x"a6",x"c4",x"7e"),
  1345 => (x"72",x"78",x"bf",x"6e"),
  1346 => (x"ed",x"e3",x"c1",x"1e"),
  1347 => (x"49",x"66",x"c8",x"48"),
  1348 => (x"20",x"4a",x"a1",x"c8"),
  1349 => (x"05",x"aa",x"71",x"41"),
  1350 => (x"51",x"10",x"87",x"f9"),
  1351 => (x"c4",x"c1",x"4a",x"26"),
  1352 => (x"cc",x"c1",x"48",x"66"),
  1353 => (x"bf",x"6e",x"78",x"f4"),
  1354 => (x"74",x"81",x"c7",x"49"),
  1355 => (x"66",x"c4",x"c1",x"51"),
  1356 => (x"c1",x"81",x"c8",x"49"),
  1357 => (x"66",x"c4",x"c1",x"51"),
  1358 => (x"c0",x"81",x"c9",x"49"),
  1359 => (x"66",x"c4",x"c1",x"51"),
  1360 => (x"c0",x"81",x"ca",x"49"),
  1361 => (x"ac",x"fb",x"c0",x"51"),
  1362 => (x"c1",x"87",x"cf",x"02"),
  1363 => (x"c8",x"1e",x"d8",x"1e"),
  1364 => (x"c8",x"49",x"bf",x"66"),
  1365 => (x"87",x"f6",x"e1",x"81"),
  1366 => (x"c8",x"c1",x"86",x"c8"),
  1367 => (x"a8",x"c0",x"48",x"66"),
  1368 => (x"c8",x"87",x"c7",x"01"),
  1369 => (x"78",x"c1",x"48",x"a6"),
  1370 => (x"c8",x"c1",x"87",x"ce"),
  1371 => (x"88",x"c1",x"48",x"66"),
  1372 => (x"c3",x"58",x"a6",x"d0"),
  1373 => (x"87",x"c2",x"e1",x"87"),
  1374 => (x"c2",x"48",x"a6",x"d8"),
  1375 => (x"02",x"9c",x"74",x"78"),
  1376 => (x"c8",x"87",x"f1",x"cc"),
  1377 => (x"cc",x"c1",x"48",x"66"),
  1378 => (x"cc",x"03",x"a8",x"66"),
  1379 => (x"a6",x"dc",x"87",x"e6"),
  1380 => (x"c4",x"78",x"c0",x"48"),
  1381 => (x"ff",x"78",x"c0",x"80"),
  1382 => (x"70",x"87",x"ca",x"df"),
  1383 => (x"48",x"66",x"d4",x"4c"),
  1384 => (x"c7",x"05",x"a8",x"dd"),
  1385 => (x"a6",x"e0",x"c0",x"87"),
  1386 => (x"78",x"66",x"d4",x"48"),
  1387 => (x"05",x"ac",x"d0",x"c1"),
  1388 => (x"ff",x"87",x"eb",x"c0"),
  1389 => (x"ff",x"87",x"ee",x"de"),
  1390 => (x"70",x"87",x"ea",x"de"),
  1391 => (x"ac",x"ec",x"c0",x"4c"),
  1392 => (x"ff",x"87",x"c6",x"05"),
  1393 => (x"70",x"87",x"f3",x"df"),
  1394 => (x"ac",x"d0",x"c1",x"4c"),
  1395 => (x"d0",x"87",x"c8",x"05"),
  1396 => (x"80",x"c1",x"48",x"66"),
  1397 => (x"c1",x"58",x"a6",x"d4"),
  1398 => (x"ff",x"02",x"ac",x"d0"),
  1399 => (x"e4",x"c0",x"87",x"d5"),
  1400 => (x"66",x"d4",x"48",x"a6"),
  1401 => (x"66",x"e0",x"c0",x"78"),
  1402 => (x"66",x"e4",x"c0",x"48"),
  1403 => (x"d5",x"ca",x"05",x"a8"),
  1404 => (x"a6",x"e8",x"c0",x"87"),
  1405 => (x"ff",x"78",x"c0",x"48"),
  1406 => (x"78",x"c0",x"80",x"dc"),
  1407 => (x"fb",x"c0",x"4d",x"74"),
  1408 => (x"db",x"c9",x"02",x"8d"),
  1409 => (x"02",x"8d",x"c9",x"87"),
  1410 => (x"8d",x"c2",x"87",x"db"),
  1411 => (x"87",x"f7",x"c1",x"02"),
  1412 => (x"c4",x"02",x"8d",x"c9"),
  1413 => (x"8d",x"c4",x"87",x"d8"),
  1414 => (x"87",x"c1",x"c1",x"02"),
  1415 => (x"c4",x"02",x"8d",x"c1"),
  1416 => (x"f5",x"c8",x"87",x"cc"),
  1417 => (x"49",x"66",x"c8",x"87"),
  1418 => (x"c4",x"c1",x"91",x"cb"),
  1419 => (x"a1",x"c4",x"81",x"66"),
  1420 => (x"71",x"7e",x"6a",x"4a"),
  1421 => (x"f9",x"e3",x"c1",x"1e"),
  1422 => (x"49",x"66",x"c4",x"48"),
  1423 => (x"20",x"4a",x"a1",x"cc"),
  1424 => (x"05",x"aa",x"71",x"41"),
  1425 => (x"10",x"87",x"f8",x"ff"),
  1426 => (x"c1",x"49",x"26",x"51"),
  1427 => (x"ff",x"79",x"d9",x"d2"),
  1428 => (x"70",x"87",x"d2",x"dc"),
  1429 => (x"48",x"a6",x"c4",x"4c"),
  1430 => (x"c3",x"c8",x"78",x"c1"),
  1431 => (x"48",x"a6",x"dc",x"87"),
  1432 => (x"ff",x"78",x"f0",x"c0"),
  1433 => (x"70",x"87",x"fe",x"db"),
  1434 => (x"ac",x"ec",x"c0",x"4c"),
  1435 => (x"87",x"c4",x"c0",x"02"),
  1436 => (x"5c",x"a6",x"e0",x"c0"),
  1437 => (x"02",x"ac",x"ec",x"c0"),
  1438 => (x"db",x"ff",x"87",x"cd"),
  1439 => (x"4c",x"70",x"87",x"e7"),
  1440 => (x"05",x"ac",x"ec",x"c0"),
  1441 => (x"c0",x"87",x"f3",x"ff"),
  1442 => (x"c0",x"02",x"ac",x"ec"),
  1443 => (x"db",x"ff",x"87",x"c4"),
  1444 => (x"1e",x"c0",x"87",x"d3"),
  1445 => (x"66",x"d0",x"1e",x"ca"),
  1446 => (x"c1",x"91",x"cb",x"49"),
  1447 => (x"71",x"48",x"66",x"cc"),
  1448 => (x"58",x"a6",x"cc",x"80"),
  1449 => (x"c4",x"48",x"66",x"c8"),
  1450 => (x"58",x"a6",x"d0",x"80"),
  1451 => (x"49",x"bf",x"66",x"cc"),
  1452 => (x"87",x"da",x"dc",x"ff"),
  1453 => (x"1e",x"de",x"1e",x"c1"),
  1454 => (x"49",x"bf",x"66",x"d4"),
  1455 => (x"87",x"ce",x"dc",x"ff"),
  1456 => (x"49",x"70",x"86",x"d0"),
  1457 => (x"c0",x"89",x"09",x"c0"),
  1458 => (x"c0",x"59",x"a6",x"f0"),
  1459 => (x"c0",x"48",x"66",x"ec"),
  1460 => (x"ee",x"c0",x"06",x"a8"),
  1461 => (x"66",x"ec",x"c0",x"87"),
  1462 => (x"03",x"a8",x"dd",x"48"),
  1463 => (x"c4",x"87",x"e4",x"c0"),
  1464 => (x"c0",x"49",x"bf",x"66"),
  1465 => (x"c0",x"81",x"66",x"ec"),
  1466 => (x"ec",x"c0",x"51",x"e0"),
  1467 => (x"81",x"c1",x"49",x"66"),
  1468 => (x"81",x"bf",x"66",x"c4"),
  1469 => (x"c0",x"51",x"c1",x"c2"),
  1470 => (x"c2",x"49",x"66",x"ec"),
  1471 => (x"bf",x"66",x"c4",x"81"),
  1472 => (x"6e",x"51",x"c0",x"81"),
  1473 => (x"f4",x"cc",x"c1",x"48"),
  1474 => (x"c8",x"49",x"6e",x"78"),
  1475 => (x"51",x"66",x"d8",x"81"),
  1476 => (x"81",x"c9",x"49",x"6e"),
  1477 => (x"6e",x"51",x"66",x"d0"),
  1478 => (x"dc",x"81",x"ca",x"49"),
  1479 => (x"66",x"d8",x"51",x"66"),
  1480 => (x"dc",x"80",x"c1",x"48"),
  1481 => (x"ec",x"48",x"58",x"a6"),
  1482 => (x"c4",x"78",x"c1",x"80"),
  1483 => (x"dc",x"ff",x"87",x"f2"),
  1484 => (x"49",x"70",x"87",x"cb"),
  1485 => (x"59",x"a6",x"f0",x"c0"),
  1486 => (x"87",x"c1",x"dc",x"ff"),
  1487 => (x"e0",x"c0",x"49",x"70"),
  1488 => (x"66",x"dc",x"59",x"a6"),
  1489 => (x"a8",x"ec",x"c0",x"48"),
  1490 => (x"87",x"ca",x"c0",x"05"),
  1491 => (x"c0",x"48",x"a6",x"dc"),
  1492 => (x"c0",x"78",x"66",x"ec"),
  1493 => (x"d8",x"ff",x"87",x"c4"),
  1494 => (x"66",x"c8",x"87",x"cb"),
  1495 => (x"c1",x"91",x"cb",x"49"),
  1496 => (x"71",x"48",x"66",x"c4"),
  1497 => (x"6e",x"7e",x"70",x"80"),
  1498 => (x"6e",x"82",x"c8",x"4a"),
  1499 => (x"c0",x"81",x"ca",x"49"),
  1500 => (x"dc",x"51",x"66",x"ec"),
  1501 => (x"81",x"c1",x"49",x"66"),
  1502 => (x"89",x"66",x"ec",x"c0"),
  1503 => (x"30",x"71",x"48",x"c1"),
  1504 => (x"89",x"c1",x"49",x"70"),
  1505 => (x"c2",x"7a",x"97",x"71"),
  1506 => (x"49",x"bf",x"e0",x"f5"),
  1507 => (x"29",x"66",x"ec",x"c0"),
  1508 => (x"48",x"4a",x"6a",x"97"),
  1509 => (x"f4",x"c0",x"98",x"71"),
  1510 => (x"49",x"6e",x"58",x"a6"),
  1511 => (x"48",x"a6",x"81",x"c4"),
  1512 => (x"e4",x"c0",x"78",x"69"),
  1513 => (x"e0",x"c0",x"48",x"66"),
  1514 => (x"c0",x"02",x"a8",x"66"),
  1515 => (x"a6",x"dc",x"87",x"c8"),
  1516 => (x"c0",x"78",x"c0",x"48"),
  1517 => (x"a6",x"dc",x"87",x"c5"),
  1518 => (x"dc",x"78",x"c1",x"48"),
  1519 => (x"e0",x"c0",x"1e",x"66"),
  1520 => (x"49",x"66",x"cc",x"1e"),
  1521 => (x"87",x"c6",x"d8",x"ff"),
  1522 => (x"4c",x"70",x"86",x"c8"),
  1523 => (x"06",x"ac",x"b7",x"c0"),
  1524 => (x"c4",x"87",x"db",x"c1"),
  1525 => (x"80",x"74",x"48",x"66"),
  1526 => (x"c0",x"58",x"a6",x"c8"),
  1527 => (x"89",x"74",x"49",x"e0"),
  1528 => (x"c1",x"4b",x"66",x"c4"),
  1529 => (x"71",x"4a",x"f6",x"e3"),
  1530 => (x"87",x"fc",x"e2",x"fe"),
  1531 => (x"c2",x"48",x"66",x"c4"),
  1532 => (x"58",x"a6",x"c8",x"80"),
  1533 => (x"48",x"66",x"e8",x"c0"),
  1534 => (x"ec",x"c0",x"80",x"c1"),
  1535 => (x"f0",x"c0",x"58",x"a6"),
  1536 => (x"81",x"c1",x"49",x"66"),
  1537 => (x"c0",x"02",x"a9",x"70"),
  1538 => (x"4d",x"c0",x"87",x"c5"),
  1539 => (x"c1",x"87",x"c2",x"c0"),
  1540 => (x"c2",x"1e",x"75",x"4d"),
  1541 => (x"e0",x"c0",x"49",x"a4"),
  1542 => (x"70",x"88",x"71",x"48"),
  1543 => (x"66",x"cc",x"1e",x"49"),
  1544 => (x"e9",x"d6",x"ff",x"49"),
  1545 => (x"c0",x"86",x"c8",x"87"),
  1546 => (x"ff",x"01",x"a8",x"b7"),
  1547 => (x"e8",x"c0",x"87",x"c6"),
  1548 => (x"d1",x"c0",x"02",x"66"),
  1549 => (x"c9",x"49",x"6e",x"87"),
  1550 => (x"66",x"e8",x"c0",x"81"),
  1551 => (x"c1",x"48",x"6e",x"51"),
  1552 => (x"c0",x"78",x"c5",x"cf"),
  1553 => (x"49",x"6e",x"87",x"cc"),
  1554 => (x"51",x"c2",x"81",x"c9"),
  1555 => (x"cf",x"c1",x"48",x"6e"),
  1556 => (x"a6",x"c4",x"78",x"f9"),
  1557 => (x"c0",x"78",x"c1",x"48"),
  1558 => (x"d5",x"ff",x"87",x"c6"),
  1559 => (x"4c",x"70",x"87",x"dc"),
  1560 => (x"c0",x"02",x"66",x"c4"),
  1561 => (x"66",x"c8",x"87",x"f5"),
  1562 => (x"a8",x"66",x"cc",x"48"),
  1563 => (x"87",x"cb",x"c0",x"04"),
  1564 => (x"c1",x"48",x"66",x"c8"),
  1565 => (x"58",x"a6",x"cc",x"80"),
  1566 => (x"cc",x"87",x"e0",x"c0"),
  1567 => (x"88",x"c1",x"48",x"66"),
  1568 => (x"c0",x"58",x"a6",x"d0"),
  1569 => (x"c6",x"c1",x"87",x"d5"),
  1570 => (x"c8",x"c0",x"05",x"ac"),
  1571 => (x"48",x"66",x"d8",x"87"),
  1572 => (x"a6",x"dc",x"80",x"c1"),
  1573 => (x"e1",x"d4",x"ff",x"58"),
  1574 => (x"d0",x"4c",x"70",x"87"),
  1575 => (x"80",x"c1",x"48",x"66"),
  1576 => (x"74",x"58",x"a6",x"d4"),
  1577 => (x"cb",x"c0",x"02",x"9c"),
  1578 => (x"48",x"66",x"c8",x"87"),
  1579 => (x"a8",x"66",x"cc",x"c1"),
  1580 => (x"87",x"da",x"f3",x"04"),
  1581 => (x"87",x"f9",x"d3",x"ff"),
  1582 => (x"c7",x"48",x"66",x"c8"),
  1583 => (x"e5",x"c0",x"03",x"a8"),
  1584 => (x"f4",x"f1",x"c2",x"87"),
  1585 => (x"c8",x"78",x"c0",x"48"),
  1586 => (x"91",x"cb",x"49",x"66"),
  1587 => (x"81",x"66",x"c4",x"c1"),
  1588 => (x"6a",x"4a",x"a1",x"c4"),
  1589 => (x"79",x"52",x"c0",x"4a"),
  1590 => (x"c1",x"48",x"66",x"c8"),
  1591 => (x"58",x"a6",x"cc",x"80"),
  1592 => (x"ff",x"04",x"a8",x"c7"),
  1593 => (x"cc",x"ff",x"87",x"db"),
  1594 => (x"f6",x"df",x"ff",x"8e"),
  1595 => (x"61",x"6f",x"4c",x"87"),
  1596 => (x"2e",x"2a",x"20",x"64"),
  1597 => (x"20",x"3a",x"00",x"20"),
  1598 => (x"50",x"49",x"44",x"00"),
  1599 => (x"69",x"77",x"53",x"20"),
  1600 => (x"65",x"68",x"63",x"74"),
  1601 => (x"73",x"1e",x"00",x"73"),
  1602 => (x"9b",x"4b",x"71",x"1e"),
  1603 => (x"c2",x"87",x"c6",x"02"),
  1604 => (x"c0",x"48",x"f0",x"f1"),
  1605 => (x"c2",x"1e",x"c7",x"78"),
  1606 => (x"49",x"bf",x"f0",x"f1"),
  1607 => (x"d7",x"e7",x"c1",x"1e"),
  1608 => (x"d8",x"f1",x"c2",x"1e"),
  1609 => (x"c9",x"ee",x"49",x"bf"),
  1610 => (x"c2",x"86",x"cc",x"87"),
  1611 => (x"49",x"bf",x"d8",x"f1"),
  1612 => (x"73",x"87",x"ea",x"e9"),
  1613 => (x"87",x"c8",x"02",x"9b"),
  1614 => (x"49",x"d7",x"e7",x"c1"),
  1615 => (x"87",x"d2",x"ed",x"c0"),
  1616 => (x"87",x"e3",x"de",x"ff"),
  1617 => (x"87",x"c9",x"c7",x"1e"),
  1618 => (x"f9",x"fe",x"49",x"c1"),
  1619 => (x"e5",x"e5",x"fe",x"87"),
  1620 => (x"02",x"98",x"70",x"87"),
  1621 => (x"ec",x"fe",x"87",x"cd"),
  1622 => (x"98",x"70",x"87",x"fe"),
  1623 => (x"c1",x"87",x"c4",x"02"),
  1624 => (x"c0",x"87",x"c2",x"4a"),
  1625 => (x"05",x"9a",x"72",x"4a"),
  1626 => (x"1e",x"c0",x"87",x"ce"),
  1627 => (x"49",x"d5",x"e6",x"c1"),
  1628 => (x"87",x"fc",x"f8",x"c0"),
  1629 => (x"87",x"fe",x"86",x"c4"),
  1630 => (x"e6",x"c1",x"1e",x"c0"),
  1631 => (x"f8",x"c0",x"49",x"e0"),
  1632 => (x"1e",x"c0",x"87",x"ee"),
  1633 => (x"87",x"c4",x"fd",x"c0"),
  1634 => (x"f8",x"c0",x"49",x"70"),
  1635 => (x"ff",x"c2",x"87",x"e2"),
  1636 => (x"26",x"8e",x"f8",x"87"),
  1637 => (x"20",x"44",x"53",x"4f"),
  1638 => (x"6c",x"69",x"61",x"66"),
  1639 => (x"00",x"2e",x"64",x"65"),
  1640 => (x"74",x"6f",x"6f",x"42"),
  1641 => (x"2e",x"67",x"6e",x"69"),
  1642 => (x"1e",x"00",x"2e",x"2e"),
  1643 => (x"48",x"f0",x"f1",x"c2"),
  1644 => (x"f1",x"c2",x"78",x"c0"),
  1645 => (x"78",x"c0",x"48",x"d8"),
  1646 => (x"c0",x"87",x"c9",x"fe"),
  1647 => (x"c0",x"87",x"ec",x"fc"),
  1648 => (x"00",x"4f",x"26",x"48"),
  1649 => (x"00",x"00",x"01",x"00"),
  1650 => (x"45",x"20",x"80",x"00"),
  1651 => (x"00",x"74",x"69",x"78"),
  1652 => (x"61",x"42",x"20",x"80"),
  1653 => (x"75",x"00",x"6b",x"63"),
  1654 => (x"84",x"00",x"00",x"13"),
  1655 => (x"00",x"00",x"00",x"2c"),
  1656 => (x"13",x"75",x"00",x"00"),
  1657 => (x"2c",x"a2",x"00",x"00"),
  1658 => (x"00",x"00",x"00",x"00"),
  1659 => (x"00",x"13",x"75",x"00"),
  1660 => (x"00",x"2c",x"c0",x"00"),
  1661 => (x"00",x"00",x"00",x"00"),
  1662 => (x"00",x"00",x"13",x"75"),
  1663 => (x"00",x"00",x"2c",x"de"),
  1664 => (x"75",x"00",x"00",x"00"),
  1665 => (x"fc",x"00",x"00",x"13"),
  1666 => (x"00",x"00",x"00",x"2c"),
  1667 => (x"13",x"75",x"00",x"00"),
  1668 => (x"2d",x"1a",x"00",x"00"),
  1669 => (x"00",x"00",x"00",x"00"),
  1670 => (x"00",x"13",x"75",x"00"),
  1671 => (x"00",x"2d",x"38",x"00"),
  1672 => (x"00",x"00",x"00",x"00"),
  1673 => (x"00",x"00",x"13",x"75"),
  1674 => (x"00",x"00",x"00",x"00"),
  1675 => (x"0a",x"00",x"00",x"00"),
  1676 => (x"00",x"00",x"00",x"14"),
  1677 => (x"00",x"00",x"00",x"00"),
  1678 => (x"fe",x"1e",x"00",x"00"),
  1679 => (x"78",x"c0",x"48",x"f0"),
  1680 => (x"09",x"79",x"09",x"cd"),
  1681 => (x"1e",x"1e",x"4f",x"26"),
  1682 => (x"7e",x"bf",x"f0",x"fe"),
  1683 => (x"4f",x"26",x"26",x"48"),
  1684 => (x"48",x"f0",x"fe",x"1e"),
  1685 => (x"4f",x"26",x"78",x"c1"),
  1686 => (x"48",x"f0",x"fe",x"1e"),
  1687 => (x"4f",x"26",x"78",x"c0"),
  1688 => (x"c0",x"4a",x"71",x"1e"),
  1689 => (x"4f",x"26",x"52",x"52"),
  1690 => (x"5c",x"5b",x"5e",x"0e"),
  1691 => (x"86",x"f4",x"0e",x"5d"),
  1692 => (x"6d",x"97",x"4d",x"71"),
  1693 => (x"4c",x"a5",x"c1",x"7e"),
  1694 => (x"c8",x"48",x"6c",x"97"),
  1695 => (x"48",x"6e",x"58",x"a6"),
  1696 => (x"05",x"a8",x"66",x"c4"),
  1697 => (x"48",x"ff",x"87",x"c5"),
  1698 => (x"ff",x"87",x"e6",x"c0"),
  1699 => (x"a5",x"c2",x"87",x"ca"),
  1700 => (x"4b",x"6c",x"97",x"49"),
  1701 => (x"97",x"4b",x"a3",x"71"),
  1702 => (x"6c",x"97",x"4b",x"6b"),
  1703 => (x"c1",x"48",x"6e",x"7e"),
  1704 => (x"58",x"a6",x"c8",x"80"),
  1705 => (x"a6",x"cc",x"98",x"c7"),
  1706 => (x"7c",x"97",x"70",x"58"),
  1707 => (x"73",x"87",x"e1",x"fe"),
  1708 => (x"26",x"8e",x"f4",x"48"),
  1709 => (x"26",x"4c",x"26",x"4d"),
  1710 => (x"0e",x"4f",x"26",x"4b"),
  1711 => (x"0e",x"5c",x"5b",x"5e"),
  1712 => (x"4c",x"71",x"86",x"f4"),
  1713 => (x"c3",x"4a",x"66",x"d8"),
  1714 => (x"a4",x"c2",x"9a",x"ff"),
  1715 => (x"49",x"6c",x"97",x"4b"),
  1716 => (x"72",x"49",x"a1",x"73"),
  1717 => (x"7e",x"6c",x"97",x"51"),
  1718 => (x"80",x"c1",x"48",x"6e"),
  1719 => (x"c7",x"58",x"a6",x"c8"),
  1720 => (x"58",x"a6",x"cc",x"98"),
  1721 => (x"8e",x"f4",x"54",x"70"),
  1722 => (x"1e",x"87",x"ca",x"ff"),
  1723 => (x"87",x"e8",x"fd",x"1e"),
  1724 => (x"49",x"4a",x"bf",x"e0"),
  1725 => (x"99",x"c0",x"e0",x"c0"),
  1726 => (x"72",x"87",x"cb",x"02"),
  1727 => (x"d6",x"f5",x"c2",x"1e"),
  1728 => (x"87",x"f7",x"fe",x"49"),
  1729 => (x"fd",x"fc",x"86",x"c4"),
  1730 => (x"fd",x"7e",x"70",x"87"),
  1731 => (x"26",x"26",x"87",x"c2"),
  1732 => (x"f5",x"c2",x"1e",x"4f"),
  1733 => (x"c7",x"fd",x"49",x"d6"),
  1734 => (x"eb",x"eb",x"c1",x"87"),
  1735 => (x"87",x"da",x"fc",x"49"),
  1736 => (x"26",x"87",x"f7",x"c3"),
  1737 => (x"5b",x"5e",x"0e",x"4f"),
  1738 => (x"71",x"0e",x"5d",x"5c"),
  1739 => (x"d6",x"f5",x"c2",x"4d"),
  1740 => (x"87",x"f4",x"fc",x"49"),
  1741 => (x"b7",x"c0",x"4b",x"70"),
  1742 => (x"c2",x"c3",x"04",x"ab"),
  1743 => (x"ab",x"f0",x"c3",x"87"),
  1744 => (x"c1",x"87",x"c9",x"05"),
  1745 => (x"c1",x"48",x"c9",x"f0"),
  1746 => (x"87",x"e3",x"c2",x"78"),
  1747 => (x"05",x"ab",x"e0",x"c3"),
  1748 => (x"f0",x"c1",x"87",x"c9"),
  1749 => (x"78",x"c1",x"48",x"cd"),
  1750 => (x"c1",x"87",x"d4",x"c2"),
  1751 => (x"02",x"bf",x"cd",x"f0"),
  1752 => (x"c0",x"c2",x"87",x"c6"),
  1753 => (x"87",x"c2",x"4c",x"a3"),
  1754 => (x"f0",x"c1",x"4c",x"73"),
  1755 => (x"c0",x"02",x"bf",x"c9"),
  1756 => (x"49",x"74",x"87",x"e0"),
  1757 => (x"91",x"29",x"b7",x"c4"),
  1758 => (x"81",x"e9",x"f1",x"c1"),
  1759 => (x"9a",x"cf",x"4a",x"74"),
  1760 => (x"48",x"c1",x"92",x"c2"),
  1761 => (x"4a",x"70",x"30",x"72"),
  1762 => (x"48",x"72",x"ba",x"ff"),
  1763 => (x"79",x"70",x"98",x"69"),
  1764 => (x"49",x"74",x"87",x"db"),
  1765 => (x"91",x"29",x"b7",x"c4"),
  1766 => (x"81",x"e9",x"f1",x"c1"),
  1767 => (x"9a",x"cf",x"4a",x"74"),
  1768 => (x"48",x"c3",x"92",x"c2"),
  1769 => (x"4a",x"70",x"30",x"72"),
  1770 => (x"70",x"b0",x"69",x"48"),
  1771 => (x"05",x"9d",x"75",x"79"),
  1772 => (x"ff",x"87",x"f0",x"c0"),
  1773 => (x"e1",x"c8",x"48",x"d0"),
  1774 => (x"48",x"d4",x"ff",x"78"),
  1775 => (x"f0",x"c1",x"78",x"c5"),
  1776 => (x"c3",x"02",x"bf",x"cd"),
  1777 => (x"78",x"e0",x"c3",x"87"),
  1778 => (x"bf",x"c9",x"f0",x"c1"),
  1779 => (x"ff",x"87",x"c6",x"02"),
  1780 => (x"f0",x"c3",x"48",x"d4"),
  1781 => (x"48",x"d4",x"ff",x"78"),
  1782 => (x"d0",x"ff",x"78",x"73"),
  1783 => (x"78",x"e1",x"c8",x"48"),
  1784 => (x"c1",x"78",x"e0",x"c0"),
  1785 => (x"c0",x"48",x"cd",x"f0"),
  1786 => (x"c9",x"f0",x"c1",x"78"),
  1787 => (x"c2",x"78",x"c0",x"48"),
  1788 => (x"f9",x"49",x"d6",x"f5"),
  1789 => (x"4b",x"70",x"87",x"f2"),
  1790 => (x"03",x"ab",x"b7",x"c0"),
  1791 => (x"c0",x"87",x"fe",x"fc"),
  1792 => (x"26",x"4d",x"26",x"48"),
  1793 => (x"26",x"4b",x"26",x"4c"),
  1794 => (x"00",x"00",x"00",x"4f"),
  1795 => (x"00",x"00",x"00",x"00"),
  1796 => (x"4a",x"71",x"1e",x"00"),
  1797 => (x"87",x"cd",x"fc",x"49"),
  1798 => (x"c0",x"1e",x"4f",x"26"),
  1799 => (x"c4",x"49",x"72",x"4a"),
  1800 => (x"e9",x"f1",x"c1",x"91"),
  1801 => (x"c1",x"79",x"c0",x"81"),
  1802 => (x"aa",x"b7",x"d0",x"82"),
  1803 => (x"26",x"87",x"ee",x"04"),
  1804 => (x"5b",x"5e",x"0e",x"4f"),
  1805 => (x"71",x"0e",x"5d",x"5c"),
  1806 => (x"87",x"dc",x"f8",x"4d"),
  1807 => (x"b7",x"c4",x"4a",x"75"),
  1808 => (x"f1",x"c1",x"92",x"2a"),
  1809 => (x"4c",x"75",x"82",x"e9"),
  1810 => (x"94",x"c2",x"9c",x"cf"),
  1811 => (x"74",x"4b",x"49",x"6a"),
  1812 => (x"c2",x"9b",x"c3",x"2b"),
  1813 => (x"70",x"30",x"74",x"48"),
  1814 => (x"74",x"bc",x"ff",x"4c"),
  1815 => (x"70",x"98",x"71",x"48"),
  1816 => (x"87",x"ec",x"f7",x"7a"),
  1817 => (x"d8",x"fe",x"48",x"73"),
  1818 => (x"00",x"00",x"00",x"87"),
  1819 => (x"00",x"00",x"00",x"00"),
  1820 => (x"00",x"00",x"00",x"00"),
  1821 => (x"00",x"00",x"00",x"00"),
  1822 => (x"00",x"00",x"00",x"00"),
  1823 => (x"00",x"00",x"00",x"00"),
  1824 => (x"00",x"00",x"00",x"00"),
  1825 => (x"00",x"00",x"00",x"00"),
  1826 => (x"00",x"00",x"00",x"00"),
  1827 => (x"00",x"00",x"00",x"00"),
  1828 => (x"00",x"00",x"00",x"00"),
  1829 => (x"00",x"00",x"00",x"00"),
  1830 => (x"00",x"00",x"00",x"00"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"00",x"00"),
  1834 => (x"d0",x"ff",x"1e",x"00"),
  1835 => (x"78",x"e1",x"c8",x"48"),
  1836 => (x"d4",x"ff",x"48",x"71"),
  1837 => (x"66",x"c4",x"78",x"08"),
  1838 => (x"08",x"d4",x"ff",x"48"),
  1839 => (x"1e",x"4f",x"26",x"78"),
  1840 => (x"66",x"c4",x"4a",x"71"),
  1841 => (x"49",x"72",x"1e",x"49"),
  1842 => (x"ff",x"87",x"de",x"ff"),
  1843 => (x"e0",x"c0",x"48",x"d0"),
  1844 => (x"4f",x"26",x"26",x"78"),
  1845 => (x"71",x"1e",x"73",x"1e"),
  1846 => (x"49",x"66",x"c8",x"4b"),
  1847 => (x"c1",x"4a",x"73",x"1e"),
  1848 => (x"ff",x"49",x"a2",x"e0"),
  1849 => (x"c4",x"26",x"87",x"d9"),
  1850 => (x"26",x"4d",x"26",x"87"),
  1851 => (x"26",x"4b",x"26",x"4c"),
  1852 => (x"d4",x"ff",x"1e",x"4f"),
  1853 => (x"7a",x"ff",x"c3",x"4a"),
  1854 => (x"c0",x"48",x"d0",x"ff"),
  1855 => (x"7a",x"de",x"78",x"e1"),
  1856 => (x"bf",x"e0",x"f5",x"c2"),
  1857 => (x"c8",x"48",x"49",x"7a"),
  1858 => (x"71",x"7a",x"70",x"28"),
  1859 => (x"70",x"28",x"d0",x"48"),
  1860 => (x"d8",x"48",x"71",x"7a"),
  1861 => (x"ff",x"7a",x"70",x"28"),
  1862 => (x"e0",x"c0",x"48",x"d0"),
  1863 => (x"0e",x"4f",x"26",x"78"),
  1864 => (x"5d",x"5c",x"5b",x"5e"),
  1865 => (x"c2",x"4c",x"71",x"0e"),
  1866 => (x"4d",x"bf",x"e0",x"f5"),
  1867 => (x"71",x"29",x"74",x"49"),
  1868 => (x"9b",x"66",x"d0",x"4b"),
  1869 => (x"66",x"d4",x"83",x"c1"),
  1870 => (x"c2",x"04",x"ab",x"b7"),
  1871 => (x"d0",x"4b",x"c0",x"87"),
  1872 => (x"31",x"74",x"49",x"66"),
  1873 => (x"99",x"75",x"b9",x"ff"),
  1874 => (x"32",x"74",x"4a",x"73"),
  1875 => (x"b0",x"71",x"48",x"72"),
  1876 => (x"58",x"e4",x"f5",x"c2"),
  1877 => (x"26",x"87",x"da",x"fe"),
  1878 => (x"26",x"4c",x"26",x"4d"),
  1879 => (x"0e",x"4f",x"26",x"4b"),
  1880 => (x"5d",x"5c",x"5b",x"5e"),
  1881 => (x"4c",x"71",x"1e",x"0e"),
  1882 => (x"4b",x"e4",x"f5",x"c2"),
  1883 => (x"f4",x"c0",x"4a",x"c0"),
  1884 => (x"c3",x"cd",x"fe",x"49"),
  1885 => (x"c2",x"1e",x"74",x"87"),
  1886 => (x"fe",x"49",x"e4",x"f5"),
  1887 => (x"c4",x"87",x"c6",x"e8"),
  1888 => (x"99",x"49",x"70",x"86"),
  1889 => (x"87",x"ea",x"c0",x"02"),
  1890 => (x"4d",x"a6",x"1e",x"c4"),
  1891 => (x"e4",x"f5",x"c2",x"1e"),
  1892 => (x"d4",x"ef",x"fe",x"49"),
  1893 => (x"70",x"86",x"c8",x"87"),
  1894 => (x"87",x"d6",x"02",x"98"),
  1895 => (x"f7",x"c1",x"4a",x"75"),
  1896 => (x"4b",x"c4",x"49",x"e8"),
  1897 => (x"87",x"c2",x"cb",x"fe"),
  1898 => (x"ca",x"02",x"98",x"70"),
  1899 => (x"c0",x"48",x"c0",x"87"),
  1900 => (x"48",x"c0",x"87",x"ed"),
  1901 => (x"c0",x"87",x"e8",x"c0"),
  1902 => (x"c4",x"c1",x"87",x"f3"),
  1903 => (x"02",x"98",x"70",x"87"),
  1904 => (x"fc",x"c0",x"87",x"c8"),
  1905 => (x"05",x"98",x"70",x"87"),
  1906 => (x"f6",x"c2",x"87",x"f8"),
  1907 => (x"cc",x"02",x"bf",x"c4"),
  1908 => (x"e0",x"f5",x"c2",x"87"),
  1909 => (x"c4",x"f6",x"c2",x"48"),
  1910 => (x"d4",x"fc",x"78",x"bf"),
  1911 => (x"26",x"48",x"c1",x"87"),
  1912 => (x"4c",x"26",x"4d",x"26"),
  1913 => (x"4f",x"26",x"4b",x"26"),
  1914 => (x"43",x"52",x"41",x"5b"),
  1915 => (x"1e",x"c0",x"1e",x"00"),
  1916 => (x"49",x"e4",x"f5",x"c2"),
  1917 => (x"87",x"cf",x"ec",x"fe"),
  1918 => (x"48",x"fc",x"f5",x"c2"),
  1919 => (x"26",x"26",x"78",x"c0"),
  1920 => (x"5b",x"5e",x"0e",x"4f"),
  1921 => (x"f4",x"0e",x"5d",x"5c"),
  1922 => (x"c2",x"7e",x"c0",x"86"),
  1923 => (x"48",x"bf",x"fc",x"f5"),
  1924 => (x"03",x"a8",x"b7",x"c3"),
  1925 => (x"f5",x"c2",x"87",x"d1"),
  1926 => (x"c1",x"48",x"bf",x"fc"),
  1927 => (x"c0",x"f6",x"c2",x"80"),
  1928 => (x"48",x"fb",x"c0",x"58"),
  1929 => (x"c2",x"87",x"d9",x"c6"),
  1930 => (x"fe",x"49",x"e4",x"f5"),
  1931 => (x"70",x"87",x"ce",x"f1"),
  1932 => (x"ac",x"b7",x"c0",x"4c"),
  1933 => (x"48",x"87",x"c4",x"03"),
  1934 => (x"c2",x"87",x"c5",x"c6"),
  1935 => (x"4a",x"bf",x"fc",x"f5"),
  1936 => (x"d8",x"02",x"8a",x"c3"),
  1937 => (x"02",x"8a",x"c1",x"87"),
  1938 => (x"8a",x"87",x"c7",x"c5"),
  1939 => (x"87",x"f2",x"c2",x"02"),
  1940 => (x"cf",x"c1",x"02",x"8a"),
  1941 => (x"c3",x"02",x"8a",x"87"),
  1942 => (x"d9",x"c5",x"87",x"de"),
  1943 => (x"c8",x"4d",x"c0",x"87"),
  1944 => (x"4a",x"75",x"5c",x"a6"),
  1945 => (x"ff",x"c1",x"92",x"c4"),
  1946 => (x"f5",x"c2",x"82",x"de"),
  1947 => (x"84",x"75",x"4c",x"f8"),
  1948 => (x"49",x"4b",x"6c",x"97"),
  1949 => (x"97",x"a3",x"c1",x"4b"),
  1950 => (x"11",x"81",x"6a",x"7c"),
  1951 => (x"58",x"a6",x"cc",x"48"),
  1952 => (x"c8",x"48",x"66",x"c4"),
  1953 => (x"c3",x"02",x"a8",x"66"),
  1954 => (x"7c",x"97",x"c0",x"87"),
  1955 => (x"c7",x"05",x"66",x"c8"),
  1956 => (x"fc",x"f5",x"c2",x"87"),
  1957 => (x"78",x"a5",x"c4",x"48"),
  1958 => (x"b7",x"c4",x"85",x"c1"),
  1959 => (x"c1",x"ff",x"04",x"ad"),
  1960 => (x"87",x"d2",x"c4",x"87"),
  1961 => (x"bf",x"c8",x"f6",x"c2"),
  1962 => (x"a8",x"b7",x"c8",x"48"),
  1963 => (x"ca",x"87",x"cb",x"01"),
  1964 => (x"87",x"c6",x"02",x"ac"),
  1965 => (x"c0",x"05",x"ac",x"cd"),
  1966 => (x"f6",x"c2",x"87",x"f3"),
  1967 => (x"c8",x"4b",x"bf",x"c8"),
  1968 => (x"d2",x"03",x"ab",x"b7"),
  1969 => (x"cc",x"f6",x"c2",x"87"),
  1970 => (x"c0",x"81",x"73",x"49"),
  1971 => (x"83",x"c1",x"51",x"e0"),
  1972 => (x"04",x"ab",x"b7",x"c8"),
  1973 => (x"c2",x"87",x"ee",x"ff"),
  1974 => (x"c1",x"48",x"d4",x"f6"),
  1975 => (x"cf",x"c1",x"50",x"d2"),
  1976 => (x"50",x"cd",x"c1",x"50"),
  1977 => (x"80",x"e4",x"50",x"c0"),
  1978 => (x"c9",x"c3",x"78",x"c3"),
  1979 => (x"c8",x"f6",x"c2",x"87"),
  1980 => (x"c1",x"48",x"49",x"bf"),
  1981 => (x"cc",x"f6",x"c2",x"80"),
  1982 => (x"a0",x"c4",x"48",x"58"),
  1983 => (x"c2",x"51",x"74",x"81"),
  1984 => (x"f0",x"c0",x"87",x"f4"),
  1985 => (x"da",x"04",x"ac",x"b7"),
  1986 => (x"b7",x"f9",x"c0",x"87"),
  1987 => (x"87",x"d3",x"01",x"ac"),
  1988 => (x"bf",x"c0",x"f6",x"c2"),
  1989 => (x"74",x"91",x"ca",x"49"),
  1990 => (x"8a",x"f0",x"c0",x"4a"),
  1991 => (x"48",x"c0",x"f6",x"c2"),
  1992 => (x"ca",x"78",x"a1",x"72"),
  1993 => (x"c6",x"c0",x"02",x"ac"),
  1994 => (x"05",x"ac",x"cd",x"87"),
  1995 => (x"c2",x"87",x"c7",x"c2"),
  1996 => (x"c3",x"48",x"fc",x"f5"),
  1997 => (x"87",x"fe",x"c1",x"78"),
  1998 => (x"ac",x"b7",x"f0",x"c0"),
  1999 => (x"c0",x"87",x"db",x"04"),
  2000 => (x"01",x"ac",x"b7",x"f9"),
  2001 => (x"c2",x"87",x"d3",x"c0"),
  2002 => (x"49",x"bf",x"c4",x"f6"),
  2003 => (x"4a",x"74",x"91",x"d0"),
  2004 => (x"c2",x"8a",x"f0",x"c0"),
  2005 => (x"72",x"48",x"c4",x"f6"),
  2006 => (x"c1",x"c1",x"78",x"a1"),
  2007 => (x"c0",x"04",x"ac",x"b7"),
  2008 => (x"c6",x"c1",x"87",x"db"),
  2009 => (x"c0",x"01",x"ac",x"b7"),
  2010 => (x"f6",x"c2",x"87",x"d3"),
  2011 => (x"d0",x"49",x"bf",x"c4"),
  2012 => (x"c0",x"4a",x"74",x"91"),
  2013 => (x"f6",x"c2",x"8a",x"f7"),
  2014 => (x"a1",x"72",x"48",x"c4"),
  2015 => (x"02",x"ac",x"ca",x"78"),
  2016 => (x"cd",x"87",x"c6",x"c0"),
  2017 => (x"ed",x"c0",x"05",x"ac"),
  2018 => (x"fc",x"f5",x"c2",x"87"),
  2019 => (x"c0",x"78",x"c3",x"48"),
  2020 => (x"e2",x"c0",x"87",x"e4"),
  2021 => (x"c6",x"c0",x"05",x"ac"),
  2022 => (x"7e",x"fb",x"c0",x"87"),
  2023 => (x"ca",x"87",x"d7",x"c0"),
  2024 => (x"c6",x"c0",x"02",x"ac"),
  2025 => (x"05",x"ac",x"cd",x"87"),
  2026 => (x"c2",x"87",x"c9",x"c0"),
  2027 => (x"c3",x"48",x"fc",x"f5"),
  2028 => (x"87",x"c2",x"c0",x"78"),
  2029 => (x"02",x"6e",x"7e",x"74"),
  2030 => (x"6e",x"87",x"d0",x"f9"),
  2031 => (x"99",x"ff",x"c3",x"48"),
  2032 => (x"db",x"f8",x"8e",x"f4"),
  2033 => (x"4e",x"4f",x"43",x"87"),
  2034 => (x"4d",x"00",x"3d",x"46"),
  2035 => (x"4e",x"00",x"44",x"4f"),
  2036 => (x"00",x"45",x"4d",x"41"),
  2037 => (x"41",x"46",x"45",x"44"),
  2038 => (x"3d",x"54",x"4c",x"55"),
  2039 => (x"1f",x"c5",x"00",x"30"),
  2040 => (x"1f",x"cb",x"00",x"00"),
  2041 => (x"1f",x"cf",x"00",x"00"),
  2042 => (x"1f",x"d4",x"00",x"00"),
  2043 => (x"ff",x"1e",x"00",x"00"),
  2044 => (x"c9",x"c8",x"48",x"d0"),
  2045 => (x"ff",x"48",x"71",x"78"),
  2046 => (x"26",x"78",x"08",x"d4"),
  2047 => (x"4a",x"71",x"1e",x"4f"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

